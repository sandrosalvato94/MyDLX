
module MUX21_31 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_30 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_29 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_28 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_27 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_26 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_25 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_24 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_23 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_22 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_21 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  AOI22_X1 U1 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U2 ( .A(S), .ZN(n1) );
  INV_X1 U3 ( .A(n2), .ZN(Y) );
endmodule


module MUX21_20 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_19 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_18 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_17 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  AOI22_X1 U1 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U2 ( .A(S), .ZN(n1) );
  INV_X1 U3 ( .A(n2), .ZN(Y) );
endmodule


module MUX21_16 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_15 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_14 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_13 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  AOI22_X1 U1 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U2 ( .A(S), .ZN(n1) );
  INV_X1 U3 ( .A(n2), .ZN(Y) );
endmodule


module MUX21_12 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_11 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_10 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_9 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  AOI22_X1 U1 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U2 ( .A(S), .ZN(n1) );
  INV_X1 U3 ( .A(n2), .ZN(Y) );
endmodule


module MUX21_8 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_7 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_6 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_5 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  AOI22_X1 U1 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U2 ( .A(S), .ZN(n1) );
  INV_X1 U3 ( .A(n2), .ZN(Y) );
endmodule


module MUX21_4 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_3 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_2 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module MUX21_1 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n2) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module FA_63 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_62 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_61 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_60 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_59 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_58 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_57 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_56 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_55 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_54 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_53 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_52 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_51 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_50 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_49 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_48 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_47 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_46 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_45 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_44 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_43 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_42 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_41 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_40 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_39 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_38 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_37 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_36 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_35 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_34 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_33 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_32 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_31 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_30 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_29 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_28 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_27 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_26 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_25 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_24 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_23 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_22 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_21 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_20 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_19 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_18 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_17 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_16 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_15 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_14 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_13 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_12 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_11 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_10 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_9 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_8 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_7 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_6 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_5 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_4 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_3 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_2 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module FA_1 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n4, n5;

  XOR2_X1 U3 ( .A(Ci), .B(n5), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n5) );
  INV_X1 U1 ( .A(n4), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n5), .B2(Ci), .ZN(n4) );
endmodule


module MUX21_GENERIC_N4_7 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_28 U_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_27 U_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_26 U_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_25 U_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_6 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_24 U_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_23 U_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_22 U_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_21 U_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_5 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_20 U_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_19 U_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_18 U_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_17 U_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_4 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_16 U_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_15 U_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_14 U_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_13 U_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_3 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_12 U_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_11 U_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_10 U_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_9 U_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_2 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_8 U_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_7 U_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_6 U_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_5 U_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module MUX21_GENERIC_N4_1 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_4 U_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_3 U_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_2 U_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_1 U_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module RCA_N4_15 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_60 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_59 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_58 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_57 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_N4_14 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_56 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_55 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_54 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_53 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_N4_13 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_52 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_51 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_50 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_49 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_N4_12 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_48 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_47 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_46 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_45 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_N4_11 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_44 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_43 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_42 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_41 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_N4_10 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_40 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_39 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_38 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_37 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_N4_9 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_36 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_35 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_34 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_33 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_N4_8 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_32 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_31 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_30 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_29 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_N4_7 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_28 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_27 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_26 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_25 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_N4_6 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_24 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_23 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_22 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_21 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_N4_5 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_20 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_19 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_18 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_17 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_N4_4 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_16 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_15 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_14 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_13 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_N4_3 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_12 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_11 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_10 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_9 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_N4_2 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_8 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_7 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_6 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_5 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module RCA_N4_1 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_4 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_3 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_2 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_1 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module CarrySelectBlock_N4_7 ( A, B, Cin, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;

  wire   [3:0] sum1;
  wire   [3:0] sum2;

  RCA_N4_14 rca1 ( .A(A), .B(B), .Ci(1'b0), .S(sum1) );
  RCA_N4_13 rca2 ( .A(A), .B(B), .Ci(1'b1), .S(sum2) );
  MUX21_GENERIC_N4_7 mux ( .A(sum1), .B(sum2), .SEL(Cin), .Y(S) );
endmodule


module CarrySelectBlock_N4_6 ( A, B, Cin, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;

  wire   [3:0] sum1;
  wire   [3:0] sum2;

  RCA_N4_12 rca1 ( .A(A), .B(B), .Ci(1'b0), .S(sum1) );
  RCA_N4_11 rca2 ( .A(A), .B(B), .Ci(1'b1), .S(sum2) );
  MUX21_GENERIC_N4_6 mux ( .A(sum1), .B(sum2), .SEL(Cin), .Y(S) );
endmodule


module CarrySelectBlock_N4_5 ( A, B, Cin, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;

  wire   [3:0] sum1;
  wire   [3:0] sum2;

  RCA_N4_10 rca1 ( .A(A), .B(B), .Ci(1'b0), .S(sum1) );
  RCA_N4_9 rca2 ( .A(A), .B(B), .Ci(1'b1), .S(sum2) );
  MUX21_GENERIC_N4_5 mux ( .A(sum1), .B(sum2), .SEL(Cin), .Y(S) );
endmodule


module CarrySelectBlock_N4_4 ( A, B, Cin, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;

  wire   [3:0] sum1;
  wire   [3:0] sum2;

  RCA_N4_8 rca1 ( .A(A), .B(B), .Ci(1'b0), .S(sum1) );
  RCA_N4_7 rca2 ( .A(A), .B(B), .Ci(1'b1), .S(sum2) );
  MUX21_GENERIC_N4_4 mux ( .A(sum1), .B(sum2), .SEL(Cin), .Y(S) );
endmodule


module CarrySelectBlock_N4_3 ( A, B, Cin, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;

  wire   [3:0] sum1;
  wire   [3:0] sum2;

  RCA_N4_6 rca1 ( .A(A), .B(B), .Ci(1'b0), .S(sum1) );
  RCA_N4_5 rca2 ( .A(A), .B(B), .Ci(1'b1), .S(sum2) );
  MUX21_GENERIC_N4_3 mux ( .A(sum1), .B(sum2), .SEL(Cin), .Y(S) );
endmodule


module CarrySelectBlock_N4_2 ( A, B, Cin, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;

  wire   [3:0] sum1;
  wire   [3:0] sum2;

  RCA_N4_4 rca1 ( .A(A), .B(B), .Ci(1'b0), .S(sum1) );
  RCA_N4_3 rca2 ( .A(A), .B(B), .Ci(1'b1), .S(sum2) );
  MUX21_GENERIC_N4_2 mux ( .A(sum1), .B(sum2), .SEL(Cin), .Y(S) );
endmodule


module CarrySelectBlock_N4_1 ( A, B, Cin, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;

  wire   [3:0] sum1;
  wire   [3:0] sum2;

  RCA_N4_2 rca1 ( .A(A), .B(B), .Ci(1'b0), .S(sum1) );
  RCA_N4_1 rca2 ( .A(A), .B(B), .Ci(1'b1), .S(sum2) );
  MUX21_GENERIC_N4_1 mux ( .A(sum1), .B(sum2), .SEL(Cin), .Y(S) );
endmodule


module GeneralPropagate_26 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_25 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_24 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_23 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_22 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_21 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  AND2_X1 U1 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
  INV_X1 U2 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U3 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
endmodule


module GeneralPropagate_20 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_19 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_18 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  AND2_X1 U1 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
  INV_X1 U2 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U3 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
endmodule


module GeneralPropagate_17 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  AND2_X1 U1 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
  INV_X1 U2 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U3 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
endmodule


module GeneralPropagate_16 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_15 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_14 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_13 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_12 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  AND2_X1 U1 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
  INV_X1 U2 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U3 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
endmodule


module GeneralPropagate_11 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_10 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_9 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_8 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_7 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_6 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  AOI21_X1 U1 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(G_ij) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_5 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  AND2_X1 U1 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
  INV_X1 U2 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U3 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
endmodule


module GeneralPropagate_4 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_3 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
  AND2_X1 U3 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
endmodule


module GeneralPropagate_2 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  AND2_X1 U1 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
  INV_X1 U2 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U3 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
endmodule


module GeneralPropagate_1 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n3;

  AND2_X1 U1 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
  INV_X1 U2 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U3 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n3) );
endmodule


module Mux_NBit_2x1_NBIT_IN40_3 ( port0, port1, sel, portY );
  input [39:0] port0;
  input [39:0] port1;
  output [39:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n43, n52, n53, n54, n55, n56,
         n57, n58, n59, n60;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;
  assign portY[32] = N34;
  assign portY[33] = N35;
  assign portY[34] = N36;
  assign portY[35] = N37;
  assign portY[36] = N38;
  assign portY[37] = N39;
  assign portY[38] = N40;
  assign portY[39] = N41;

  BUF_X2 U1 ( .A(n1), .Z(n9) );
  CLKBUF_X1 U2 ( .A(n9), .Z(n11) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n1) );
  BUF_X2 U4 ( .A(sel), .Z(n2) );
  BUF_X1 U5 ( .A(n2), .Z(n7) );
  INV_X2 U6 ( .A(n2), .ZN(n5) );
  INV_X1 U7 ( .A(n2), .ZN(n4) );
  INV_X1 U8 ( .A(n2), .ZN(n3) );
  BUF_X1 U9 ( .A(n2), .Z(n10) );
  BUF_X1 U10 ( .A(n2), .Z(n8) );
  INV_X1 U11 ( .A(n34), .ZN(N30) );
  INV_X1 U12 ( .A(n32), .ZN(N29) );
  INV_X1 U13 ( .A(n30), .ZN(N27) );
  INV_X1 U14 ( .A(n35), .ZN(N31) );
  INV_X1 U15 ( .A(n54), .ZN(N40) );
  INV_X1 U16 ( .A(n55), .ZN(N41) );
  AOI22_X1 U17 ( .A1(port0[39]), .A2(n3), .B1(port1[39]), .B2(n7), .ZN(n55) );
  INV_X1 U18 ( .A(n29), .ZN(N26) );
  AOI22_X1 U19 ( .A1(port0[29]), .A2(n6), .B1(port1[29]), .B2(n8), .ZN(n35) );
  AOI22_X1 U20 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n8), .ZN(n34) );
  AOI22_X1 U21 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n9), .ZN(n32) );
  AOI22_X1 U22 ( .A1(port0[25]), .A2(n3), .B1(port1[25]), .B2(n9), .ZN(n30) );
  AOI22_X1 U23 ( .A1(port0[35]), .A2(n4), .B1(port1[35]), .B2(n10), .ZN(n41)
         );
  INV_X1 U24 ( .A(n31), .ZN(N28) );
  AOI22_X1 U25 ( .A1(port0[33]), .A2(n4), .B1(port1[33]), .B2(n1), .ZN(n39) );
  AOI22_X1 U26 ( .A1(port0[37]), .A2(n6), .B1(port1[37]), .B2(n7), .ZN(n52) );
  AOI22_X1 U27 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n10), .ZN(n29)
         );
  INV_X1 U28 ( .A(n27), .ZN(N24) );
  INV_X1 U29 ( .A(n25), .ZN(N22) );
  INV_X1 U30 ( .A(n26), .ZN(N23) );
  INV_X1 U31 ( .A(n20), .ZN(N18) );
  INV_X1 U32 ( .A(n23), .ZN(N20) );
  INV_X1 U33 ( .A(n21), .ZN(N19) );
  INV_X1 U34 ( .A(n19), .ZN(N17) );
  INV_X1 U35 ( .A(n18), .ZN(N16) );
  INV_X1 U36 ( .A(n14), .ZN(N12) );
  INV_X1 U37 ( .A(n17), .ZN(N15) );
  INV_X1 U38 ( .A(n16), .ZN(N14) );
  INV_X1 U39 ( .A(n15), .ZN(N13) );
  INV_X1 U40 ( .A(n28), .ZN(N25) );
  INV_X1 U41 ( .A(n24), .ZN(N21) );
  INV_X1 U42 ( .A(n13), .ZN(N11) );
  INV_X1 U43 ( .A(n22), .ZN(N2) );
  INV_X1 U44 ( .A(n12), .ZN(N10) );
  INV_X1 U45 ( .A(n56), .ZN(N5) );
  INV_X1 U46 ( .A(n53), .ZN(N4) );
  INV_X1 U47 ( .A(n33), .ZN(N3) );
  INV_X1 U48 ( .A(n60), .ZN(N9) );
  INV_X1 U49 ( .A(n59), .ZN(N8) );
  INV_X1 U50 ( .A(n58), .ZN(N7) );
  INV_X1 U51 ( .A(n57), .ZN(N6) );
  AOI22_X1 U52 ( .A1(port0[26]), .A2(n6), .B1(port1[26]), .B2(n9), .ZN(n31) );
  AOI22_X1 U53 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n10), .ZN(n28)
         );
  AOI22_X1 U54 ( .A1(port0[16]), .A2(n5), .B1(port1[16]), .B2(n11), .ZN(n20)
         );
  AOI22_X1 U55 ( .A1(port0[22]), .A2(n6), .B1(port1[22]), .B2(n10), .ZN(n27)
         );
  AOI22_X1 U56 ( .A1(port0[21]), .A2(n3), .B1(port1[21]), .B2(n9), .ZN(n26) );
  AOI22_X1 U57 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n11), .ZN(n25)
         );
  AOI22_X1 U58 ( .A1(port0[18]), .A2(n6), .B1(port1[18]), .B2(n11), .ZN(n23)
         );
  AOI22_X1 U59 ( .A1(port0[15]), .A2(n5), .B1(port1[15]), .B2(n11), .ZN(n19)
         );
  AOI22_X1 U60 ( .A1(port0[17]), .A2(n3), .B1(port1[17]), .B2(n11), .ZN(n21)
         );
  AOI22_X1 U61 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n11), .ZN(n24)
         );
  AOI22_X1 U62 ( .A1(port0[14]), .A2(n6), .B1(port1[14]), .B2(n11), .ZN(n18)
         );
  AOI22_X1 U63 ( .A1(port0[9]), .A2(n5), .B1(port1[9]), .B2(n11), .ZN(n13) );
  AOI22_X1 U64 ( .A1(port0[10]), .A2(n6), .B1(port1[10]), .B2(n11), .ZN(n14)
         );
  AOI22_X1 U65 ( .A1(port0[13]), .A2(n3), .B1(port1[13]), .B2(n11), .ZN(n17)
         );
  AOI22_X1 U66 ( .A1(port0[12]), .A2(n5), .B1(port1[12]), .B2(n11), .ZN(n16)
         );
  AOI22_X1 U67 ( .A1(port0[11]), .A2(n6), .B1(port1[11]), .B2(n11), .ZN(n15)
         );
  AOI22_X1 U68 ( .A1(port0[1]), .A2(n3), .B1(port1[1]), .B2(n9), .ZN(n33) );
  AOI22_X1 U69 ( .A1(port0[0]), .A2(n6), .B1(port1[0]), .B2(n11), .ZN(n22) );
  AOI22_X1 U70 ( .A1(port0[8]), .A2(n3), .B1(port1[8]), .B2(n11), .ZN(n12) );
  AOI22_X1 U71 ( .A1(port0[3]), .A2(n6), .B1(port1[3]), .B2(n7), .ZN(n56) );
  AOI22_X1 U72 ( .A1(port0[2]), .A2(n3), .B1(port1[2]), .B2(n11), .ZN(n53) );
  AOI22_X1 U73 ( .A1(port0[7]), .A2(n3), .B1(n11), .B2(port1[7]), .ZN(n60) );
  AOI22_X1 U74 ( .A1(port0[6]), .A2(n5), .B1(port1[6]), .B2(n11), .ZN(n59) );
  AOI22_X1 U75 ( .A1(port0[5]), .A2(n6), .B1(port1[5]), .B2(n7), .ZN(n58) );
  AOI22_X1 U76 ( .A1(port0[4]), .A2(n3), .B1(port1[4]), .B2(n11), .ZN(n57) );
  AOI22_X1 U77 ( .A1(port0[34]), .A2(n4), .B1(port1[34]), .B2(n1), .ZN(n40) );
  AOI22_X1 U78 ( .A1(port0[36]), .A2(n5), .B1(port1[36]), .B2(n7), .ZN(n43) );
  AOI22_X1 U79 ( .A1(port0[31]), .A2(n4), .B1(port1[31]), .B2(n8), .ZN(n37) );
  AOI22_X1 U80 ( .A1(port0[38]), .A2(n3), .B1(port1[38]), .B2(n9), .ZN(n54) );
  AOI22_X1 U81 ( .A1(port0[32]), .A2(n4), .B1(port1[32]), .B2(n1), .ZN(n38) );
  INV_X1 U82 ( .A(n36), .ZN(N32) );
  INV_X1 U83 ( .A(n52), .ZN(N39) );
  INV_X1 U84 ( .A(n43), .ZN(N38) );
  INV_X1 U85 ( .A(n38), .ZN(N34) );
  AOI22_X1 U86 ( .A1(port0[30]), .A2(n4), .B1(port1[30]), .B2(n8), .ZN(n36) );
  INV_X1 U87 ( .A(n40), .ZN(N36) );
  INV_X1 U88 ( .A(n41), .ZN(N37) );
  INV_X1 U89 ( .A(n39), .ZN(N35) );
  INV_X1 U90 ( .A(n37), .ZN(N33) );
  INV_X1 U91 ( .A(n2), .ZN(n6) );
endmodule


module Mux_NBit_2x1_NBIT_IN40_2 ( port0, port1, sel, portY );
  input [39:0] port0;
  input [39:0] port1;
  output [39:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, n1, n2, n3, n4,
         n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n43, n52, n53, n54, n55, n56,
         n57, n58, n59, n60;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;
  assign portY[32] = N34;
  assign portY[33] = N35;
  assign portY[34] = N36;
  assign portY[35] = N37;
  assign portY[36] = N38;
  assign portY[37] = N39;
  assign portY[38] = N40;
  assign portY[39] = N41;

  BUF_X1 U1 ( .A(sel), .Z(n2) );
  BUF_X1 U2 ( .A(n1), .Z(n10) );
  INV_X1 U3 ( .A(n6), .ZN(n3) );
  BUF_X1 U4 ( .A(n1), .Z(n11) );
  BUF_X1 U5 ( .A(n1), .Z(n9) );
  BUF_X1 U6 ( .A(sel), .Z(n8) );
  BUF_X1 U7 ( .A(n2), .Z(n7) );
  INV_X1 U8 ( .A(n55), .ZN(N41) );
  CLKBUF_X1 U9 ( .A(n10), .Z(n6) );
  INV_X1 U10 ( .A(n34), .ZN(N30) );
  INV_X1 U11 ( .A(n32), .ZN(N29) );
  AOI22_X1 U12 ( .A1(port0[27]), .A2(n4), .B1(port1[27]), .B2(n10), .ZN(n32)
         );
  INV_X1 U13 ( .A(n30), .ZN(N27) );
  AOI22_X1 U14 ( .A1(port0[25]), .A2(n4), .B1(port1[25]), .B2(n10), .ZN(n30)
         );
  INV_X1 U15 ( .A(n35), .ZN(N31) );
  INV_X1 U16 ( .A(n54), .ZN(N40) );
  BUF_X1 U17 ( .A(sel), .Z(n1) );
  INV_X1 U18 ( .A(n29), .ZN(N26) );
  AOI22_X1 U19 ( .A1(port0[24]), .A2(n4), .B1(port1[24]), .B2(n11), .ZN(n29)
         );
  INV_X1 U20 ( .A(n31), .ZN(N28) );
  AOI22_X1 U21 ( .A1(port0[26]), .A2(n4), .B1(port1[26]), .B2(n10), .ZN(n31)
         );
  INV_X1 U22 ( .A(n27), .ZN(N24) );
  AOI22_X1 U23 ( .A1(port0[22]), .A2(n4), .B1(port1[22]), .B2(n11), .ZN(n27)
         );
  INV_X1 U24 ( .A(n25), .ZN(N22) );
  AOI22_X1 U25 ( .A1(port0[20]), .A2(n4), .B1(port1[20]), .B2(n6), .ZN(n25) );
  INV_X1 U26 ( .A(n26), .ZN(N23) );
  AOI22_X1 U27 ( .A1(port0[21]), .A2(n4), .B1(port1[21]), .B2(n6), .ZN(n26) );
  INV_X1 U28 ( .A(n20), .ZN(N18) );
  AOI22_X1 U29 ( .A1(port0[16]), .A2(n3), .B1(port1[16]), .B2(n6), .ZN(n20) );
  INV_X1 U30 ( .A(n23), .ZN(N20) );
  AOI22_X1 U31 ( .A1(port0[18]), .A2(n3), .B1(port1[18]), .B2(n6), .ZN(n23) );
  INV_X1 U32 ( .A(n21), .ZN(N19) );
  AOI22_X1 U33 ( .A1(port0[17]), .A2(n3), .B1(port1[17]), .B2(n6), .ZN(n21) );
  INV_X1 U34 ( .A(n19), .ZN(N17) );
  AOI22_X1 U35 ( .A1(port0[15]), .A2(n3), .B1(port1[15]), .B2(n6), .ZN(n19) );
  INV_X1 U36 ( .A(n18), .ZN(N16) );
  AOI22_X1 U37 ( .A1(port0[14]), .A2(n3), .B1(port1[14]), .B2(n6), .ZN(n18) );
  INV_X1 U38 ( .A(n14), .ZN(N12) );
  AOI22_X1 U39 ( .A1(port0[10]), .A2(n3), .B1(port1[10]), .B2(n6), .ZN(n14) );
  INV_X1 U40 ( .A(n17), .ZN(N15) );
  AOI22_X1 U41 ( .A1(port0[13]), .A2(n3), .B1(port1[13]), .B2(n6), .ZN(n17) );
  INV_X1 U42 ( .A(n16), .ZN(N14) );
  AOI22_X1 U43 ( .A1(port0[12]), .A2(n3), .B1(port1[12]), .B2(n6), .ZN(n16) );
  INV_X1 U44 ( .A(n15), .ZN(N13) );
  AOI22_X1 U45 ( .A1(port0[11]), .A2(n3), .B1(port1[11]), .B2(n6), .ZN(n15) );
  INV_X1 U46 ( .A(n28), .ZN(N25) );
  AOI22_X1 U47 ( .A1(port0[23]), .A2(n4), .B1(port1[23]), .B2(n11), .ZN(n28)
         );
  INV_X1 U48 ( .A(n24), .ZN(N21) );
  AOI22_X1 U49 ( .A1(port0[19]), .A2(n4), .B1(port1[19]), .B2(n6), .ZN(n24) );
  INV_X1 U50 ( .A(n13), .ZN(N11) );
  AOI22_X1 U51 ( .A1(port0[9]), .A2(n3), .B1(port1[9]), .B2(n6), .ZN(n13) );
  INV_X1 U52 ( .A(n22), .ZN(N2) );
  AOI22_X1 U53 ( .A1(port0[0]), .A2(n3), .B1(port1[0]), .B2(n6), .ZN(n22) );
  INV_X1 U54 ( .A(n12), .ZN(N10) );
  AOI22_X1 U55 ( .A1(port0[8]), .A2(n3), .B1(port1[8]), .B2(n6), .ZN(n12) );
  INV_X1 U56 ( .A(n56), .ZN(N5) );
  INV_X1 U57 ( .A(n53), .ZN(N4) );
  INV_X1 U58 ( .A(n33), .ZN(N3) );
  AOI22_X1 U59 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n10), .ZN(n33) );
  INV_X1 U60 ( .A(n60), .ZN(N9) );
  AOI22_X1 U61 ( .A1(port0[7]), .A2(n3), .B1(n6), .B2(port1[7]), .ZN(n60) );
  INV_X1 U62 ( .A(n59), .ZN(N8) );
  AOI22_X1 U63 ( .A1(port0[6]), .A2(n3), .B1(port1[6]), .B2(n6), .ZN(n59) );
  INV_X1 U64 ( .A(n58), .ZN(N7) );
  AOI22_X1 U65 ( .A1(port0[5]), .A2(n3), .B1(port1[5]), .B2(n6), .ZN(n58) );
  INV_X1 U66 ( .A(n57), .ZN(N6) );
  AOI22_X1 U67 ( .A1(port0[4]), .A2(n3), .B1(port1[4]), .B2(n6), .ZN(n57) );
  AOI22_X1 U68 ( .A1(port0[28]), .A2(n4), .B1(port1[28]), .B2(n9), .ZN(n34) );
  AOI22_X1 U69 ( .A1(port0[29]), .A2(n4), .B1(port1[29]), .B2(n9), .ZN(n35) );
  AOI22_X1 U70 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(n7), .ZN(n53) );
  AOI22_X1 U71 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n56) );
  AOI22_X1 U72 ( .A1(port0[39]), .A2(n5), .B1(port1[39]), .B2(n7), .ZN(n55) );
  AOI22_X1 U73 ( .A1(port0[38]), .A2(n5), .B1(port1[38]), .B2(n7), .ZN(n54) );
  AOI22_X1 U74 ( .A1(port0[37]), .A2(n5), .B1(port1[37]), .B2(n7), .ZN(n52) );
  AOI22_X1 U75 ( .A1(port0[34]), .A2(n5), .B1(port1[34]), .B2(n8), .ZN(n40) );
  AOI22_X1 U76 ( .A1(port0[32]), .A2(n5), .B1(port1[32]), .B2(n8), .ZN(n38) );
  AOI22_X1 U77 ( .A1(port0[36]), .A2(n5), .B1(port1[36]), .B2(n8), .ZN(n43) );
  AOI22_X1 U78 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n9), .ZN(n36) );
  AOI22_X1 U79 ( .A1(port0[35]), .A2(n5), .B1(port1[35]), .B2(n11), .ZN(n41)
         );
  AOI22_X1 U80 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n9), .ZN(n37) );
  INV_X1 U81 ( .A(n52), .ZN(N39) );
  INV_X1 U82 ( .A(n43), .ZN(N38) );
  INV_X1 U83 ( .A(n36), .ZN(N32) );
  INV_X1 U84 ( .A(n38), .ZN(N34) );
  INV_X1 U85 ( .A(n39), .ZN(N35) );
  INV_X1 U86 ( .A(n40), .ZN(N36) );
  INV_X1 U87 ( .A(n41), .ZN(N37) );
  AOI22_X1 U88 ( .A1(port0[33]), .A2(n5), .B1(port1[33]), .B2(n8), .ZN(n39) );
  INV_X1 U89 ( .A(n37), .ZN(N33) );
  INV_X2 U90 ( .A(n2), .ZN(n4) );
  INV_X2 U91 ( .A(n2), .ZN(n5) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_20 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  CLKBUF_X1 U1 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n1) );
  INV_X1 U4 ( .A(n8), .ZN(N5) );
  AOI22_X1 U5 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  INV_X1 U6 ( .A(n7), .ZN(N4) );
  AOI22_X1 U7 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  AOI22_X1 U8 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  INV_X1 U9 ( .A(n6), .ZN(N3) );
  AOI22_X1 U10 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  INV_X1 U11 ( .A(n5), .ZN(N2) );
  AOI22_X1 U12 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  INV_X1 U13 ( .A(n14), .ZN(N9) );
  AOI22_X1 U14 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  INV_X1 U15 ( .A(n13), .ZN(N8) );
  INV_X1 U16 ( .A(n11), .ZN(N7) );
  AOI22_X1 U17 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  INV_X1 U18 ( .A(n9), .ZN(N6) );
  AOI22_X1 U19 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_19 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  CLKBUF_X1 U1 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n1) );
  INV_X1 U4 ( .A(n14), .ZN(N9) );
  AOI22_X1 U5 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  INV_X1 U6 ( .A(n13), .ZN(N8) );
  AOI22_X1 U7 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  INV_X1 U8 ( .A(n6), .ZN(N3) );
  AOI22_X1 U9 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  INV_X1 U10 ( .A(n7), .ZN(N4) );
  AOI22_X1 U11 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  INV_X1 U12 ( .A(n11), .ZN(N7) );
  AOI22_X1 U13 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  INV_X1 U14 ( .A(n9), .ZN(N6) );
  AOI22_X1 U15 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  INV_X1 U16 ( .A(n8), .ZN(N5) );
  AOI22_X1 U17 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  INV_X1 U18 ( .A(n5), .ZN(N2) );
  AOI22_X1 U19 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_18 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  CLKBUF_X1 U1 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n1) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n3) );
  AOI22_X1 U4 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  AOI22_X1 U5 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  AOI22_X1 U6 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  AOI22_X1 U7 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  AOI22_X1 U8 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  INV_X1 U9 ( .A(n14), .ZN(N9) );
  INV_X1 U10 ( .A(n5), .ZN(N2) );
  INV_X1 U11 ( .A(n13), .ZN(N8) );
  INV_X1 U12 ( .A(n11), .ZN(N7) );
  INV_X1 U13 ( .A(n9), .ZN(N6) );
  AOI22_X1 U14 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  INV_X1 U15 ( .A(n7), .ZN(N4) );
  AOI22_X1 U16 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  INV_X1 U17 ( .A(n6), .ZN(N3) );
  AOI22_X1 U18 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  INV_X1 U19 ( .A(n8), .ZN(N5) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_17 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  CLKBUF_X1 U1 ( .A(sel), .Z(n2) );
  BUF_X1 U2 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n1) );
  AOI22_X1 U4 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  AOI22_X1 U5 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  INV_X1 U6 ( .A(n8), .ZN(N5) );
  AOI22_X1 U7 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  INV_X1 U8 ( .A(n7), .ZN(N4) );
  AOI22_X1 U9 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  INV_X1 U10 ( .A(n6), .ZN(N3) );
  AOI22_X1 U11 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  INV_X1 U12 ( .A(n5), .ZN(N2) );
  AOI22_X1 U13 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  INV_X1 U14 ( .A(n14), .ZN(N9) );
  INV_X1 U15 ( .A(n11), .ZN(N7) );
  INV_X1 U16 ( .A(n9), .ZN(N6) );
  INV_X1 U17 ( .A(n13), .ZN(N8) );
  AOI22_X1 U18 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  AOI22_X1 U19 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_16 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  CLKBUF_X1 U1 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n1) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n2) );
  INV_X1 U4 ( .A(n14), .ZN(N9) );
  INV_X1 U5 ( .A(n6), .ZN(N3) );
  INV_X1 U6 ( .A(n11), .ZN(N7) );
  INV_X1 U7 ( .A(n13), .ZN(N8) );
  INV_X1 U8 ( .A(n8), .ZN(N5) );
  INV_X1 U9 ( .A(n7), .ZN(N4) );
  INV_X1 U10 ( .A(n9), .ZN(N6) );
  INV_X1 U11 ( .A(n5), .ZN(N2) );
  AOI22_X1 U12 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  AOI22_X1 U13 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  AOI22_X1 U14 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  AOI22_X1 U15 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  AOI22_X1 U16 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  AOI22_X1 U17 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  AOI22_X1 U19 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_15 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  CLKBUF_X1 U1 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n1) );
  INV_X1 U4 ( .A(n8), .ZN(N5) );
  INV_X1 U5 ( .A(n7), .ZN(N4) );
  AOI22_X1 U6 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  AOI22_X1 U7 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  AOI22_X1 U8 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  AOI22_X1 U9 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  AOI22_X1 U10 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  AOI22_X1 U11 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  AOI22_X1 U12 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  INV_X1 U13 ( .A(n6), .ZN(N3) );
  INV_X1 U14 ( .A(n5), .ZN(N2) );
  INV_X1 U15 ( .A(n14), .ZN(N9) );
  INV_X1 U16 ( .A(n13), .ZN(N8) );
  AOI22_X1 U17 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  INV_X1 U18 ( .A(n11), .ZN(N7) );
  INV_X1 U19 ( .A(n9), .ZN(N6) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_14 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  CLKBUF_X1 U1 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n1) );
  INV_X1 U4 ( .A(n14), .ZN(N9) );
  INV_X1 U5 ( .A(n13), .ZN(N8) );
  INV_X1 U6 ( .A(n6), .ZN(N3) );
  INV_X1 U7 ( .A(n7), .ZN(N4) );
  INV_X1 U8 ( .A(n11), .ZN(N7) );
  INV_X1 U9 ( .A(n9), .ZN(N6) );
  INV_X1 U10 ( .A(n8), .ZN(N5) );
  INV_X1 U11 ( .A(n5), .ZN(N2) );
  AOI22_X1 U12 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  AOI22_X1 U13 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  AOI22_X1 U14 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  AOI22_X1 U15 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  AOI22_X1 U16 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  AOI22_X1 U17 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  AOI22_X1 U19 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_13 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  CLKBUF_X1 U1 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n1) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n3) );
  AOI22_X1 U4 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  AOI22_X1 U5 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  AOI22_X1 U6 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  INV_X1 U7 ( .A(n14), .ZN(N9) );
  INV_X1 U8 ( .A(n5), .ZN(N2) );
  AOI22_X1 U9 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  INV_X1 U10 ( .A(n13), .ZN(N8) );
  INV_X1 U11 ( .A(n11), .ZN(N7) );
  AOI22_X1 U12 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  INV_X1 U13 ( .A(n9), .ZN(N6) );
  INV_X1 U14 ( .A(n7), .ZN(N4) );
  INV_X1 U15 ( .A(n6), .ZN(N3) );
  INV_X1 U16 ( .A(n8), .ZN(N5) );
  AOI22_X1 U17 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  AOI22_X1 U18 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  AOI22_X1 U19 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_12 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  BUF_X1 U1 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n1) );
  INV_X1 U4 ( .A(n8), .ZN(N5) );
  INV_X1 U5 ( .A(n7), .ZN(N4) );
  INV_X1 U6 ( .A(n6), .ZN(N3) );
  INV_X1 U7 ( .A(n5), .ZN(N2) );
  INV_X1 U8 ( .A(n11), .ZN(N7) );
  INV_X1 U9 ( .A(n9), .ZN(N6) );
  INV_X1 U10 ( .A(n14), .ZN(N9) );
  INV_X1 U11 ( .A(n13), .ZN(N8) );
  AOI22_X1 U12 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  AOI22_X1 U13 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  AOI22_X1 U14 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  AOI22_X1 U15 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  AOI22_X1 U16 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  AOI22_X1 U17 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  AOI22_X1 U19 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_11 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  BUF_X1 U1 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n1) );
  INV_X1 U4 ( .A(n14), .ZN(N9) );
  INV_X1 U5 ( .A(n13), .ZN(N8) );
  INV_X1 U6 ( .A(n7), .ZN(N4) );
  INV_X1 U7 ( .A(n11), .ZN(N7) );
  INV_X1 U8 ( .A(n5), .ZN(N2) );
  INV_X1 U9 ( .A(n8), .ZN(N5) );
  INV_X1 U10 ( .A(n9), .ZN(N6) );
  AOI22_X1 U11 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  AOI22_X1 U12 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  AOI22_X1 U13 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  AOI22_X1 U14 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  AOI22_X1 U15 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  INV_X1 U16 ( .A(n6), .ZN(N3) );
  AOI22_X1 U17 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  AOI22_X1 U19 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_10 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  CLKBUF_X1 U1 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n1) );
  AOI22_X1 U4 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  AOI22_X1 U5 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  AOI22_X1 U6 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  AOI22_X1 U7 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  AOI22_X1 U8 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  AOI22_X1 U9 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  INV_X1 U10 ( .A(n6), .ZN(N3) );
  AOI22_X1 U11 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  INV_X1 U12 ( .A(n5), .ZN(N2) );
  INV_X1 U13 ( .A(n8), .ZN(N5) );
  INV_X1 U14 ( .A(n7), .ZN(N4) );
  INV_X1 U15 ( .A(n14), .ZN(N9) );
  INV_X1 U16 ( .A(n13), .ZN(N8) );
  INV_X1 U17 ( .A(n11), .ZN(N7) );
  INV_X1 U18 ( .A(n9), .ZN(N6) );
  AOI22_X1 U19 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_9 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  CLKBUF_X1 U1 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n1) );
  AOI22_X1 U4 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  INV_X1 U5 ( .A(n14), .ZN(N9) );
  INV_X1 U6 ( .A(n13), .ZN(N8) );
  INV_X1 U7 ( .A(n6), .ZN(N3) );
  AOI22_X1 U8 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  INV_X1 U9 ( .A(n7), .ZN(N4) );
  AOI22_X1 U10 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  INV_X1 U11 ( .A(n11), .ZN(N7) );
  AOI22_X1 U12 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  INV_X1 U13 ( .A(n9), .ZN(N6) );
  INV_X1 U14 ( .A(n8), .ZN(N5) );
  AOI22_X1 U15 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  INV_X1 U16 ( .A(n5), .ZN(N2) );
  AOI22_X1 U17 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  AOI22_X1 U18 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  AOI22_X1 U19 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_8 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  CLKBUF_X1 U1 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n1) );
  INV_X1 U4 ( .A(n14), .ZN(N9) );
  INV_X1 U5 ( .A(n5), .ZN(N2) );
  INV_X1 U6 ( .A(n13), .ZN(N8) );
  INV_X1 U7 ( .A(n11), .ZN(N7) );
  INV_X1 U8 ( .A(n9), .ZN(N6) );
  INV_X1 U9 ( .A(n7), .ZN(N4) );
  INV_X1 U10 ( .A(n6), .ZN(N3) );
  INV_X1 U11 ( .A(n8), .ZN(N5) );
  AOI22_X1 U12 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  AOI22_X1 U13 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  AOI22_X1 U14 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  AOI22_X1 U15 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  AOI22_X1 U16 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  AOI22_X1 U17 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  AOI22_X1 U19 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_7 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  BUF_X1 U1 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n1) );
  INV_X1 U4 ( .A(n11), .ZN(N7) );
  INV_X1 U5 ( .A(n9), .ZN(N6) );
  INV_X1 U6 ( .A(n8), .ZN(N5) );
  INV_X1 U7 ( .A(n6), .ZN(N3) );
  INV_X1 U8 ( .A(n5), .ZN(N2) );
  INV_X1 U9 ( .A(n7), .ZN(N4) );
  INV_X1 U10 ( .A(n13), .ZN(N8) );
  INV_X1 U11 ( .A(n14), .ZN(N9) );
  AOI22_X1 U12 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  AOI22_X1 U13 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  AOI22_X1 U14 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  AOI22_X1 U15 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  AOI22_X1 U16 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  AOI22_X1 U17 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  AOI22_X1 U19 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_6 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  BUF_X1 U1 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n1) );
  INV_X1 U4 ( .A(n14), .ZN(N9) );
  INV_X1 U5 ( .A(n5), .ZN(N2) );
  INV_X1 U6 ( .A(n9), .ZN(N6) );
  INV_X1 U7 ( .A(n8), .ZN(N5) );
  INV_X1 U8 ( .A(n7), .ZN(N4) );
  INV_X1 U9 ( .A(n6), .ZN(N3) );
  INV_X1 U10 ( .A(n11), .ZN(N7) );
  INV_X1 U11 ( .A(n13), .ZN(N8) );
  AOI22_X1 U12 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  AOI22_X1 U13 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  AOI22_X1 U14 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  AOI22_X1 U15 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  AOI22_X1 U16 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  AOI22_X1 U17 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  AOI22_X1 U19 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_5 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  CLKBUF_X1 U1 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n1) );
  AOI22_X1 U4 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  AOI22_X1 U5 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  INV_X1 U6 ( .A(n6), .ZN(N3) );
  INV_X1 U7 ( .A(n5), .ZN(N2) );
  AOI22_X1 U8 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  INV_X1 U9 ( .A(n8), .ZN(N5) );
  AOI22_X1 U10 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  INV_X1 U11 ( .A(n7), .ZN(N4) );
  AOI22_X1 U12 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  INV_X1 U13 ( .A(n14), .ZN(N9) );
  INV_X1 U14 ( .A(n13), .ZN(N8) );
  INV_X1 U15 ( .A(n11), .ZN(N7) );
  AOI22_X1 U16 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  INV_X1 U17 ( .A(n9), .ZN(N6) );
  AOI22_X1 U18 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  AOI22_X1 U19 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_4 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  CLKBUF_X1 U1 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n1) );
  INV_X1 U4 ( .A(n14), .ZN(N9) );
  INV_X1 U5 ( .A(n13), .ZN(N8) );
  INV_X1 U6 ( .A(n6), .ZN(N3) );
  INV_X1 U7 ( .A(n7), .ZN(N4) );
  INV_X1 U8 ( .A(n11), .ZN(N7) );
  INV_X1 U9 ( .A(n9), .ZN(N6) );
  INV_X1 U10 ( .A(n8), .ZN(N5) );
  INV_X1 U11 ( .A(n5), .ZN(N2) );
  AOI22_X1 U12 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  AOI22_X1 U13 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  AOI22_X1 U14 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  AOI22_X1 U15 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  AOI22_X1 U16 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  AOI22_X1 U17 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  AOI22_X1 U19 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_3 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  CLKBUF_X1 U1 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n1) );
  INV_X1 U4 ( .A(n14), .ZN(N9) );
  INV_X1 U5 ( .A(n5), .ZN(N2) );
  INV_X1 U6 ( .A(n13), .ZN(N8) );
  INV_X1 U7 ( .A(n11), .ZN(N7) );
  INV_X1 U8 ( .A(n9), .ZN(N6) );
  INV_X1 U9 ( .A(n7), .ZN(N4) );
  INV_X1 U10 ( .A(n6), .ZN(N3) );
  INV_X1 U11 ( .A(n8), .ZN(N5) );
  AOI22_X1 U12 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  AOI22_X1 U13 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  AOI22_X1 U14 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  AOI22_X1 U15 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  AOI22_X1 U16 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  AOI22_X1 U17 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  AOI22_X1 U19 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_2 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  BUF_X1 U1 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n1) );
  INV_X1 U4 ( .A(n11), .ZN(N7) );
  INV_X1 U5 ( .A(n9), .ZN(N6) );
  INV_X1 U6 ( .A(n8), .ZN(N5) );
  INV_X1 U7 ( .A(n6), .ZN(N3) );
  INV_X1 U8 ( .A(n5), .ZN(N2) );
  INV_X1 U9 ( .A(n7), .ZN(N4) );
  INV_X1 U10 ( .A(n14), .ZN(N9) );
  AOI22_X1 U11 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  AOI22_X1 U12 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  AOI22_X1 U13 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  AOI22_X1 U14 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  AOI22_X1 U15 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  INV_X1 U16 ( .A(n13), .ZN(N8) );
  AOI22_X1 U17 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  AOI22_X1 U19 ( .A1(port0[7]), .A2(n4), .B1(port1[7]), .B2(n3), .ZN(n14) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_1 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n11, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  CLKBUF_X1 U1 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n1) );
  CLKBUF_X1 U3 ( .A(sel), .Z(n2) );
  INV_X1 U4 ( .A(n14), .ZN(N9) );
  INV_X1 U5 ( .A(n9), .ZN(N6) );
  INV_X1 U6 ( .A(n8), .ZN(N5) );
  INV_X1 U7 ( .A(n6), .ZN(N3) );
  INV_X1 U8 ( .A(n11), .ZN(N7) );
  INV_X1 U9 ( .A(n13), .ZN(N8) );
  INV_X1 U10 ( .A(n7), .ZN(N4) );
  INV_X1 U11 ( .A(n5), .ZN(N2) );
  AOI22_X1 U12 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n2), .ZN(n6) );
  AOI22_X1 U13 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n2), .ZN(n11) );
  AOI22_X1 U14 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n2), .ZN(n9) );
  AOI22_X1 U15 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n3), .ZN(n13) );
  AOI22_X1 U16 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n1), .ZN(n5) );
  AOI22_X1 U17 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n1), .ZN(n7) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n1), .ZN(n8) );
  AOI22_X1 U19 ( .A1(port0[7]), .A2(n4), .B1(n3), .B2(port1[7]), .ZN(n14) );
  INV_X1 U20 ( .A(n3), .ZN(n4) );
endmodule


module PG_cell_92 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_91 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_90 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_89 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_88 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_87 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_86 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_85 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_84 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_83 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_82 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_81 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_80 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_79 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_78 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_77 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_76 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_75 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_74 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_73 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_72 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_71 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_70 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_69 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_68 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_67 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_66 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_65 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_64 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_63 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_62 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_61 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_60 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_59 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_58 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_57 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_56 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_55 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_54 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_53 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_52 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_51 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_50 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_49 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_48 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_47 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_46 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_45 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_44 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_43 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_42 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_41 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_40 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_39 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_38 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_37 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_36 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_35 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_34 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_33 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_32 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_31 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_30 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_29 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_28 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_27 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_26 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_25 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_24 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_23 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_22 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_21 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_20 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_19 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_18 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_17 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_16 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_15 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_14 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_13 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_12 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_11 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_10 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_9 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_8 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_7 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_6 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_5 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_4 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_3 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_2 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module PG_cell_1 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module GeneralGenerate_11 ( G_ik, P_ik, G_km1_j, G_ij );
  input G_ik, P_ik, G_km1_j;
  output G_ij;
  wire   n3;

  AOI21_X1 U1 ( .B1(P_ik), .B2(G_km1_j), .A(G_ik), .ZN(n3) );
  INV_X1 U2 ( .A(n3), .ZN(G_ij) );
endmodule


module GeneralGenerate_10 ( G_ik, P_ik, G_km1_j, G_ij );
  input G_ik, P_ik, G_km1_j;
  output G_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_km1_j), .A(G_ik), .ZN(n3) );
endmodule


module GeneralGenerate_9 ( G_ik, P_ik, G_km1_j, G_ij );
  input G_ik, P_ik, G_km1_j;
  output G_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_km1_j), .A(G_ik), .ZN(n3) );
endmodule


module GeneralGenerate_8 ( G_ik, P_ik, G_km1_j, G_ij );
  input G_ik, P_ik, G_km1_j;
  output G_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_km1_j), .A(G_ik), .ZN(n3) );
endmodule


module GeneralGenerate_7 ( G_ik, P_ik, G_km1_j, G_ij );
  input G_ik, P_ik, G_km1_j;
  output G_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_km1_j), .A(G_ik), .ZN(n3) );
endmodule


module GeneralGenerate_6 ( G_ik, P_ik, G_km1_j, G_ij );
  input G_ik, P_ik, G_km1_j;
  output G_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_km1_j), .A(G_ik), .ZN(n3) );
endmodule


module GeneralGenerate_5 ( G_ik, P_ik, G_km1_j, G_ij );
  input G_ik, P_ik, G_km1_j;
  output G_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_km1_j), .A(G_ik), .ZN(n3) );
endmodule


module GeneralGenerate_4 ( G_ik, P_ik, G_km1_j, G_ij );
  input G_ik, P_ik, G_km1_j;
  output G_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_km1_j), .A(G_ik), .ZN(n3) );
endmodule


module GeneralGenerate_3 ( G_ik, P_ik, G_km1_j, G_ij );
  input G_ik, P_ik, G_km1_j;
  output G_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_km1_j), .A(G_ik), .ZN(n3) );
endmodule


module GeneralGenerate_2 ( G_ik, P_ik, G_km1_j, G_ij );
  input G_ik, P_ik, G_km1_j;
  output G_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_km1_j), .A(G_ik), .ZN(n3) );
endmodule


module GeneralGenerate_1 ( G_ik, P_ik, G_km1_j, G_ij );
  input G_ik, P_ik, G_km1_j;
  output G_ij;
  wire   n3;

  INV_X1 U1 ( .A(n3), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_km1_j), .A(G_ik), .ZN(n3) );
endmodule


module t_ff_rst0_63 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_62 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_61 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_60 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_59 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_58 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_57 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_56 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_55 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_54 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_53 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_52 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_51 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_50 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_49 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_48 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_47 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_46 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_45 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_44 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_43 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_42 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_41 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_40 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_39 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_38 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_37 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_36 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_35 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_34 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_33 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_32 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_31 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_30 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_29 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_28 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_27 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_26 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_25 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_24 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_23 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_22 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_21 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_20 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_19 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_18 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_17 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_16 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_15 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_14 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_13 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_12 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_11 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_10 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_9 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_8 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_7 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_6 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_5 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_4 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_3 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_2 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_1 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_31 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_30 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_29 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_28 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_27 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_26 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_25 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_24 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_23 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_22 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_21 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_20 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_19 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_18 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_17 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_16 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_15 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_14 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_13 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_12 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_11 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_10 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_9 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_8 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_7 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_6 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_5 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_4 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_3 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_2 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst1_1 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN6_1 ( port0, port1, sel, portY );
  input [5:0] port0;
  input [5:0] port1;
  output [5:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, n1, n2, n3, n4, n5, n6, n7;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;

  INV_X1 U1 ( .A(sel), .ZN(n6) );
  INV_X1 U2 ( .A(n7), .ZN(N7) );
  AOI22_X1 U3 ( .A1(port0[5]), .A2(n6), .B1(sel), .B2(port1[5]), .ZN(n7) );
  INV_X1 U4 ( .A(n1), .ZN(N2) );
  AOI22_X1 U5 ( .A1(port0[0]), .A2(n6), .B1(port1[0]), .B2(sel), .ZN(n1) );
  INV_X1 U6 ( .A(n2), .ZN(N3) );
  AOI22_X1 U7 ( .A1(port0[1]), .A2(n6), .B1(port1[1]), .B2(sel), .ZN(n2) );
  INV_X1 U8 ( .A(n3), .ZN(N4) );
  AOI22_X1 U9 ( .A1(port0[2]), .A2(n6), .B1(port1[2]), .B2(sel), .ZN(n3) );
  INV_X1 U10 ( .A(n4), .ZN(N5) );
  AOI22_X1 U11 ( .A1(port0[3]), .A2(n6), .B1(port1[3]), .B2(sel), .ZN(n4) );
  INV_X1 U12 ( .A(n5), .ZN(N6) );
  AOI22_X1 U13 ( .A1(port0[4]), .A2(n6), .B1(port1[4]), .B2(sel), .ZN(n5) );
endmodule


module Mux_NBit_2x1_NBIT_IN10_1 ( port0, port1, sel, portY );
  input [9:0] port0;
  input [9:0] port1;
  output [9:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, n1, n2, n3, n4, n5, n6, n7,
         n8, n9, n10, n11;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;

  INV_X1 U1 ( .A(sel), .ZN(n10) );
  INV_X1 U2 ( .A(n7), .ZN(N6) );
  AOI22_X1 U3 ( .A1(port0[4]), .A2(n10), .B1(port1[4]), .B2(sel), .ZN(n7) );
  INV_X1 U4 ( .A(n8), .ZN(N7) );
  AOI22_X1 U5 ( .A1(port0[5]), .A2(n10), .B1(port1[5]), .B2(sel), .ZN(n8) );
  INV_X1 U6 ( .A(n3), .ZN(N2) );
  AOI22_X1 U7 ( .A1(port0[0]), .A2(n10), .B1(port1[0]), .B2(sel), .ZN(n3) );
  INV_X1 U8 ( .A(n4), .ZN(N3) );
  AOI22_X1 U9 ( .A1(port0[1]), .A2(n10), .B1(port1[1]), .B2(sel), .ZN(n4) );
  INV_X1 U10 ( .A(n5), .ZN(N4) );
  AOI22_X1 U11 ( .A1(port0[2]), .A2(n10), .B1(port1[2]), .B2(sel), .ZN(n5) );
  INV_X1 U12 ( .A(n6), .ZN(N5) );
  AOI22_X1 U13 ( .A1(port0[3]), .A2(n10), .B1(port1[3]), .B2(sel), .ZN(n6) );
  INV_X1 U14 ( .A(n11), .ZN(N9) );
  AOI22_X1 U15 ( .A1(port0[7]), .A2(n10), .B1(sel), .B2(port1[7]), .ZN(n11) );
  INV_X1 U16 ( .A(n2), .ZN(N11) );
  AOI22_X1 U17 ( .A1(port0[9]), .A2(n10), .B1(port1[9]), .B2(sel), .ZN(n2) );
  INV_X1 U18 ( .A(n9), .ZN(N8) );
  AOI22_X1 U19 ( .A1(port0[6]), .A2(n10), .B1(port1[6]), .B2(sel), .ZN(n9) );
  INV_X1 U20 ( .A(n1), .ZN(N10) );
  AOI22_X1 U21 ( .A1(port0[8]), .A2(n10), .B1(port1[8]), .B2(sel), .ZN(n1) );
endmodule


module Enable_Interface_NBIT_DATA5_1 ( EI_datain, EI_enable, EI_dataout );
  input [4:0] EI_datain;
  output [4:0] EI_dataout;
  input EI_enable;


  AND2_X1 U1 ( .A1(EI_datain[0]), .A2(EI_enable), .ZN(EI_dataout[0]) );
  AND2_X1 U2 ( .A1(EI_datain[1]), .A2(EI_enable), .ZN(EI_dataout[1]) );
  AND2_X1 U3 ( .A1(EI_datain[2]), .A2(EI_enable), .ZN(EI_dataout[2]) );
  AND2_X1 U4 ( .A1(EI_datain[3]), .A2(EI_enable), .ZN(EI_dataout[3]) );
  AND2_X1 U5 ( .A1(EI_enable), .A2(EI_datain[4]), .ZN(EI_dataout[4]) );
endmodule


module Sum_Network_N32_1 ( G, P, S );
  input [31:0] G;
  input [31:0] P;
  output [31:0] S;


  XOR2_X1 U1 ( .A(P[9]), .B(G[9]), .Z(S[9]) );
  XOR2_X1 U2 ( .A(P[8]), .B(G[8]), .Z(S[8]) );
  XOR2_X1 U3 ( .A(P[7]), .B(G[7]), .Z(S[7]) );
  XOR2_X1 U4 ( .A(P[6]), .B(G[6]), .Z(S[6]) );
  XOR2_X1 U5 ( .A(P[5]), .B(G[5]), .Z(S[5]) );
  XOR2_X1 U6 ( .A(P[4]), .B(G[4]), .Z(S[4]) );
  XOR2_X1 U7 ( .A(P[3]), .B(G[3]), .Z(S[3]) );
  XOR2_X1 U8 ( .A(G[31]), .B(P[31]), .Z(S[31]) );
  XOR2_X1 U9 ( .A(P[30]), .B(G[30]), .Z(S[30]) );
  XOR2_X1 U10 ( .A(P[2]), .B(G[2]), .Z(S[2]) );
  XOR2_X1 U11 ( .A(P[29]), .B(G[29]), .Z(S[29]) );
  XOR2_X1 U12 ( .A(P[28]), .B(G[28]), .Z(S[28]) );
  XOR2_X1 U13 ( .A(P[27]), .B(G[27]), .Z(S[27]) );
  XOR2_X1 U14 ( .A(P[26]), .B(G[26]), .Z(S[26]) );
  XOR2_X1 U15 ( .A(P[25]), .B(G[25]), .Z(S[25]) );
  XOR2_X1 U16 ( .A(P[24]), .B(G[24]), .Z(S[24]) );
  XOR2_X1 U17 ( .A(P[23]), .B(G[23]), .Z(S[23]) );
  XOR2_X1 U18 ( .A(P[22]), .B(G[22]), .Z(S[22]) );
  XOR2_X1 U19 ( .A(P[21]), .B(G[21]), .Z(S[21]) );
  XOR2_X1 U20 ( .A(P[20]), .B(G[20]), .Z(S[20]) );
  XOR2_X1 U21 ( .A(P[1]), .B(G[1]), .Z(S[1]) );
  XOR2_X1 U22 ( .A(P[19]), .B(G[19]), .Z(S[19]) );
  XOR2_X1 U23 ( .A(P[18]), .B(G[18]), .Z(S[18]) );
  XOR2_X1 U24 ( .A(P[17]), .B(G[17]), .Z(S[17]) );
  XOR2_X1 U25 ( .A(P[16]), .B(G[16]), .Z(S[16]) );
  XOR2_X1 U26 ( .A(P[15]), .B(G[15]), .Z(S[15]) );
  XOR2_X1 U27 ( .A(P[14]), .B(G[14]), .Z(S[14]) );
  XOR2_X1 U28 ( .A(P[13]), .B(G[13]), .Z(S[13]) );
  XOR2_X1 U29 ( .A(P[12]), .B(G[12]), .Z(S[12]) );
  XOR2_X1 U30 ( .A(P[11]), .B(G[11]), .Z(S[11]) );
  XOR2_X1 U31 ( .A(P[10]), .B(G[10]), .Z(S[10]) );
  XOR2_X1 U32 ( .A(P[0]), .B(G[0]), .Z(S[0]) );
endmodule


module Carry_Network_N32_1 ( G, P, Cin, Cout, Gout, Pout );
  input [31:0] G;
  input [31:0] P;
  output [31:0] Gout;
  output [31:0] Pout;
  input Cin;
  output Cout;
  wire   Cin, n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n74, n75, n77, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113;
  assign Gout[0] = Cin;
  assign Pout[31] = P[31];
  assign Pout[30] = P[30];
  assign Pout[29] = P[29];
  assign Pout[28] = P[28];
  assign Pout[27] = P[27];
  assign Pout[26] = P[26];
  assign Pout[25] = P[25];
  assign Pout[24] = P[24];
  assign Pout[23] = P[23];
  assign Pout[22] = P[22];
  assign Pout[21] = P[21];
  assign Pout[20] = P[20];
  assign Pout[19] = P[19];
  assign Pout[18] = P[18];
  assign Pout[17] = P[17];
  assign Pout[16] = P[16];
  assign Pout[15] = P[15];
  assign Pout[14] = P[14];
  assign Pout[13] = P[13];
  assign Pout[12] = P[12];
  assign Pout[11] = P[11];
  assign Pout[10] = P[10];
  assign Pout[9] = P[9];
  assign Pout[8] = P[8];
  assign Pout[7] = P[7];
  assign Pout[6] = P[6];
  assign Pout[5] = P[5];
  assign Pout[4] = P[4];
  assign Pout[3] = P[3];
  assign Pout[2] = P[2];
  assign Pout[1] = P[1];
  assign Pout[0] = P[0];

  CLKBUF_X1 U1 ( .A(n124), .Z(Gout[1]) );
  INV_X1 U2 ( .A(G[6]), .ZN(n83) );
  INV_X1 U3 ( .A(G[30]), .ZN(n80) );
  CLKBUF_X1 U4 ( .A(n122), .Z(Gout[3]) );
  CLKBUF_X1 U5 ( .A(n117), .Z(Gout[10]) );
  CLKBUF_X1 U6 ( .A(n116), .Z(Gout[11]) );
  CLKBUF_X1 U7 ( .A(n115), .Z(Gout[12]) );
  CLKBUF_X1 U8 ( .A(n114), .Z(Gout[13]) );
  CLKBUF_X1 U9 ( .A(n119), .Z(Gout[8]) );
  CLKBUF_X1 U10 ( .A(n123), .Z(Gout[2]) );
  CLKBUF_X1 U11 ( .A(n121), .Z(Gout[4]) );
  CLKBUF_X1 U12 ( .A(n118), .Z(Gout[9]) );
  CLKBUF_X1 U13 ( .A(n120), .Z(Gout[5]) );
  CLKBUF_X1 U14 ( .A(Gout[31]), .Z(n74) );
  AOI21_X1 U15 ( .B1(P[5]), .B2(Gout[5]), .A(G[5]), .ZN(n75) );
  CLKBUF_X1 U16 ( .A(n81), .Z(Gout[7]) );
  AOI21_X1 U17 ( .B1(P[29]), .B2(Gout[29]), .A(G[29]), .ZN(n77) );
  INV_X1 U18 ( .A(P[30]), .ZN(n79) );
  OAI21_X1 U19 ( .B1(n79), .B2(n112), .A(n80), .ZN(Gout[31]) );
  INV_X1 U20 ( .A(P[6]), .ZN(n82) );
  OAI21_X1 U21 ( .B1(n89), .B2(n82), .A(n83), .ZN(n81) );
  INV_X1 U22 ( .A(n113), .ZN(Cout) );
  INV_X1 U23 ( .A(n101), .ZN(Gout[19]) );
  AOI21_X1 U24 ( .B1(P[18]), .B2(Gout[18]), .A(G[18]), .ZN(n101) );
  INV_X1 U25 ( .A(n104), .ZN(Gout[22]) );
  AOI21_X1 U26 ( .B1(P[21]), .B2(Gout[21]), .A(G[21]), .ZN(n104) );
  INV_X1 U27 ( .A(n105), .ZN(Gout[23]) );
  AOI21_X1 U28 ( .B1(P[22]), .B2(Gout[22]), .A(G[22]), .ZN(n105) );
  INV_X1 U29 ( .A(n106), .ZN(Gout[24]) );
  AOI21_X1 U30 ( .B1(P[23]), .B2(Gout[23]), .A(G[23]), .ZN(n106) );
  INV_X1 U31 ( .A(n100), .ZN(Gout[18]) );
  AOI21_X1 U32 ( .B1(P[17]), .B2(Gout[17]), .A(G[17]), .ZN(n100) );
  INV_X1 U33 ( .A(n109), .ZN(Gout[27]) );
  AOI21_X1 U34 ( .B1(P[26]), .B2(Gout[26]), .A(G[26]), .ZN(n109) );
  INV_X1 U35 ( .A(n110), .ZN(Gout[28]) );
  AOI21_X1 U36 ( .B1(P[27]), .B2(Gout[27]), .A(G[27]), .ZN(n110) );
  INV_X1 U37 ( .A(n111), .ZN(Gout[29]) );
  AOI21_X1 U38 ( .B1(P[28]), .B2(Gout[28]), .A(G[28]), .ZN(n111) );
  INV_X1 U39 ( .A(n99), .ZN(Gout[17]) );
  AOI21_X1 U40 ( .B1(P[16]), .B2(Gout[16]), .A(G[16]), .ZN(n99) );
  INV_X1 U41 ( .A(n96), .ZN(Gout[14]) );
  AOI21_X1 U42 ( .B1(n114), .B2(P[13]), .A(G[13]), .ZN(n96) );
  INV_X1 U43 ( .A(n95), .ZN(n114) );
  AOI21_X1 U44 ( .B1(n115), .B2(P[12]), .A(G[12]), .ZN(n95) );
  INV_X1 U45 ( .A(n94), .ZN(n115) );
  AOI21_X1 U46 ( .B1(n116), .B2(P[11]), .A(G[11]), .ZN(n94) );
  AOI21_X1 U47 ( .B1(n121), .B2(P[4]), .A(G[4]), .ZN(n88) );
  AOI21_X1 U48 ( .B1(P[19]), .B2(Gout[19]), .A(G[19]), .ZN(n102) );
  AOI21_X1 U49 ( .B1(P[24]), .B2(Gout[24]), .A(G[24]), .ZN(n107) );
  AOI21_X1 U50 ( .B1(P[29]), .B2(Gout[29]), .A(G[29]), .ZN(n112) );
  AOI21_X1 U51 ( .B1(P[14]), .B2(Gout[14]), .A(G[14]), .ZN(n97) );
  AOI21_X1 U52 ( .B1(n118), .B2(P[9]), .A(G[9]), .ZN(n92) );
  INV_X1 U53 ( .A(n103), .ZN(Gout[21]) );
  INV_X1 U54 ( .A(n108), .ZN(Gout[26]) );
  INV_X1 U55 ( .A(n98), .ZN(Gout[16]) );
  INV_X1 U56 ( .A(n93), .ZN(n116) );
  INV_X1 U57 ( .A(n75), .ZN(Gout[6]) );
  INV_X1 U58 ( .A(n91), .ZN(n118) );
  AOI21_X1 U59 ( .B1(n119), .B2(P[8]), .A(G[8]), .ZN(n91) );
  INV_X1 U60 ( .A(n90), .ZN(n119) );
  AOI21_X1 U61 ( .B1(n81), .B2(P[7]), .A(G[7]), .ZN(n90) );
  INV_X1 U62 ( .A(n87), .ZN(n121) );
  AOI21_X1 U63 ( .B1(n122), .B2(P[3]), .A(G[3]), .ZN(n87) );
  INV_X1 U64 ( .A(n86), .ZN(n122) );
  AOI21_X1 U65 ( .B1(n123), .B2(P[2]), .A(G[2]), .ZN(n86) );
  INV_X1 U66 ( .A(n85), .ZN(n123) );
  AOI21_X1 U67 ( .B1(n124), .B2(P[1]), .A(G[1]), .ZN(n85) );
  AOI21_X1 U68 ( .B1(P[31]), .B2(n74), .A(G[31]), .ZN(n113) );
  INV_X1 U69 ( .A(n84), .ZN(n124) );
  INV_X1 U70 ( .A(n77), .ZN(Gout[30]) );
  AOI21_X1 U71 ( .B1(P[25]), .B2(Gout[25]), .A(G[25]), .ZN(n108) );
  INV_X1 U72 ( .A(n107), .ZN(Gout[25]) );
  AOI21_X1 U73 ( .B1(P[20]), .B2(Gout[20]), .A(G[20]), .ZN(n103) );
  INV_X1 U74 ( .A(n102), .ZN(Gout[20]) );
  AOI21_X1 U75 ( .B1(P[15]), .B2(Gout[15]), .A(G[15]), .ZN(n98) );
  INV_X1 U76 ( .A(n97), .ZN(Gout[15]) );
  AOI21_X1 U77 ( .B1(n117), .B2(P[10]), .A(G[10]), .ZN(n93) );
  INV_X1 U78 ( .A(n92), .ZN(n117) );
  AOI21_X1 U79 ( .B1(n120), .B2(P[5]), .A(G[5]), .ZN(n89) );
  INV_X1 U80 ( .A(n88), .ZN(n120) );
  AOI21_X1 U81 ( .B1(P[0]), .B2(Cin), .A(G[0]), .ZN(n84) );
endmodule


module PG_network_N32_2 ( A, B, c_in, G, P );
  input [31:0] A;
  input [31:0] B;
  output [31:0] G;
  output [31:0] P;
  input c_in;
  wire   tmp1, tmp2, n1;
  assign P[0] = 1'b0;

  GeneralGenerate_11 G_cell_0_0 ( .G_ik(tmp1), .P_ik(tmp2), .G_km1_j(c_in), 
        .G_ij(G[0]) );
  PG_cell_62 PG_cell_i_1 ( .A(A[1]), .B(B[1]), .p(P[1]), .g(G[1]) );
  PG_cell_61 PG_cell_i_2 ( .A(A[2]), .B(B[2]), .p(P[2]), .g(G[2]) );
  PG_cell_60 PG_cell_i_3 ( .A(A[3]), .B(B[3]), .p(P[3]), .g(G[3]) );
  PG_cell_59 PG_cell_i_4 ( .A(A[4]), .B(B[4]), .p(P[4]), .g(G[4]) );
  PG_cell_58 PG_cell_i_5 ( .A(A[5]), .B(B[5]), .p(P[5]), .g(G[5]) );
  PG_cell_57 PG_cell_i_6 ( .A(A[6]), .B(B[6]), .p(P[6]), .g(G[6]) );
  PG_cell_56 PG_cell_i_7 ( .A(A[7]), .B(B[7]), .p(P[7]), .g(G[7]) );
  PG_cell_55 PG_cell_i_8 ( .A(A[8]), .B(B[8]), .p(P[8]), .g(G[8]) );
  PG_cell_54 PG_cell_i_9 ( .A(A[9]), .B(B[9]), .p(P[9]), .g(G[9]) );
  PG_cell_53 PG_cell_i_10 ( .A(A[10]), .B(B[10]), .p(P[10]), .g(G[10]) );
  PG_cell_52 PG_cell_i_11 ( .A(A[11]), .B(B[11]), .p(P[11]), .g(G[11]) );
  PG_cell_51 PG_cell_i_12 ( .A(A[12]), .B(B[12]), .p(P[12]), .g(G[12]) );
  PG_cell_50 PG_cell_i_13 ( .A(A[13]), .B(B[13]), .p(P[13]), .g(G[13]) );
  PG_cell_49 PG_cell_i_14 ( .A(A[14]), .B(B[14]), .p(P[14]), .g(G[14]) );
  PG_cell_48 PG_cell_i_15 ( .A(A[15]), .B(B[15]), .p(P[15]), .g(G[15]) );
  PG_cell_47 PG_cell_i_16 ( .A(A[16]), .B(B[16]), .p(P[16]), .g(G[16]) );
  PG_cell_46 PG_cell_i_17 ( .A(A[17]), .B(B[17]), .p(P[17]), .g(G[17]) );
  PG_cell_45 PG_cell_i_18 ( .A(A[18]), .B(B[18]), .p(P[18]), .g(G[18]) );
  PG_cell_44 PG_cell_i_19 ( .A(A[19]), .B(B[19]), .p(P[19]), .g(G[19]) );
  PG_cell_43 PG_cell_i_20 ( .A(A[20]), .B(B[20]), .p(P[20]), .g(G[20]) );
  PG_cell_42 PG_cell_i_21 ( .A(A[21]), .B(B[21]), .p(P[21]), .g(G[21]) );
  PG_cell_41 PG_cell_i_22 ( .A(A[22]), .B(B[22]), .p(P[22]), .g(G[22]) );
  PG_cell_40 PG_cell_i_23 ( .A(A[23]), .B(B[23]), .p(P[23]), .g(G[23]) );
  PG_cell_39 PG_cell_i_24 ( .A(A[24]), .B(B[24]), .p(P[24]), .g(G[24]) );
  PG_cell_38 PG_cell_i_25 ( .A(A[25]), .B(B[25]), .p(P[25]), .g(G[25]) );
  PG_cell_37 PG_cell_i_26 ( .A(A[26]), .B(B[26]), .p(P[26]), .g(G[26]) );
  PG_cell_36 PG_cell_i_27 ( .A(A[27]), .B(B[27]), .p(P[27]), .g(G[27]) );
  PG_cell_35 PG_cell_i_28 ( .A(A[28]), .B(B[28]), .p(P[28]), .g(G[28]) );
  PG_cell_34 PG_cell_i_29 ( .A(A[29]), .B(B[29]), .p(P[29]), .g(G[29]) );
  PG_cell_33 PG_cell_i_30 ( .A(A[30]), .B(B[30]), .p(P[30]), .g(G[30]) );
  PG_cell_32 PG_cell_i_31 ( .A(A[31]), .B(B[31]), .p(P[31]), .g(G[31]) );
  INV_X1 U2 ( .A(B[0]), .ZN(n1) );
  XNOR2_X1 U3 ( .A(A[0]), .B(n1), .ZN(tmp2) );
  AND2_X1 U4 ( .A1(A[0]), .A2(B[0]), .ZN(tmp1) );
endmodule


module PG_network_N32_1 ( A, B, c_in, G, P );
  input [31:0] A;
  input [31:0] B;
  output [31:0] G;
  output [31:0] P;
  input c_in;
  wire   tmp1, tmp2;
  assign P[0] = 1'b0;

  XOR2_X1 U3 ( .A(B[0]), .B(A[0]), .Z(tmp2) );
  GeneralGenerate_1 G_cell_0_0 ( .G_ik(tmp1), .P_ik(tmp2), .G_km1_j(c_in), 
        .G_ij(G[0]) );
  PG_cell_31 PG_cell_i_1 ( .A(A[1]), .B(B[1]), .p(P[1]), .g(G[1]) );
  PG_cell_30 PG_cell_i_2 ( .A(A[2]), .B(B[2]), .p(P[2]), .g(G[2]) );
  PG_cell_29 PG_cell_i_3 ( .A(A[3]), .B(B[3]), .p(P[3]), .g(G[3]) );
  PG_cell_28 PG_cell_i_4 ( .A(A[4]), .B(B[4]), .p(P[4]), .g(G[4]) );
  PG_cell_27 PG_cell_i_5 ( .A(A[5]), .B(B[5]), .p(P[5]), .g(G[5]) );
  PG_cell_26 PG_cell_i_6 ( .A(A[6]), .B(B[6]), .p(P[6]), .g(G[6]) );
  PG_cell_25 PG_cell_i_7 ( .A(A[7]), .B(B[7]), .p(P[7]), .g(G[7]) );
  PG_cell_24 PG_cell_i_8 ( .A(A[8]), .B(B[8]), .p(P[8]), .g(G[8]) );
  PG_cell_23 PG_cell_i_9 ( .A(A[9]), .B(B[9]), .p(P[9]), .g(G[9]) );
  PG_cell_22 PG_cell_i_10 ( .A(A[10]), .B(B[10]), .p(P[10]), .g(G[10]) );
  PG_cell_21 PG_cell_i_11 ( .A(A[11]), .B(B[11]), .p(P[11]), .g(G[11]) );
  PG_cell_20 PG_cell_i_12 ( .A(A[12]), .B(B[12]), .p(P[12]), .g(G[12]) );
  PG_cell_19 PG_cell_i_13 ( .A(A[13]), .B(B[13]), .p(P[13]), .g(G[13]) );
  PG_cell_18 PG_cell_i_14 ( .A(A[14]), .B(B[14]), .p(P[14]), .g(G[14]) );
  PG_cell_17 PG_cell_i_15 ( .A(A[15]), .B(B[15]), .p(P[15]), .g(G[15]) );
  PG_cell_16 PG_cell_i_16 ( .A(A[16]), .B(B[16]), .p(P[16]), .g(G[16]) );
  PG_cell_15 PG_cell_i_17 ( .A(A[17]), .B(B[17]), .p(P[17]), .g(G[17]) );
  PG_cell_14 PG_cell_i_18 ( .A(A[18]), .B(B[18]), .p(P[18]), .g(G[18]) );
  PG_cell_13 PG_cell_i_19 ( .A(A[19]), .B(B[19]), .p(P[19]), .g(G[19]) );
  PG_cell_12 PG_cell_i_20 ( .A(A[20]), .B(B[20]), .p(P[20]), .g(G[20]) );
  PG_cell_11 PG_cell_i_21 ( .A(A[21]), .B(B[21]), .p(P[21]), .g(G[21]) );
  PG_cell_10 PG_cell_i_22 ( .A(A[22]), .B(B[22]), .p(P[22]), .g(G[22]) );
  PG_cell_9 PG_cell_i_23 ( .A(A[23]), .B(B[23]), .p(P[23]), .g(G[23]) );
  PG_cell_8 PG_cell_i_24 ( .A(A[24]), .B(B[24]), .p(P[24]), .g(G[24]) );
  PG_cell_7 PG_cell_i_25 ( .A(A[25]), .B(B[25]), .p(P[25]), .g(G[25]) );
  PG_cell_6 PG_cell_i_26 ( .A(A[26]), .B(B[26]), .p(P[26]), .g(G[26]) );
  PG_cell_5 PG_cell_i_27 ( .A(A[27]), .B(B[27]), .p(P[27]), .g(G[27]) );
  PG_cell_4 PG_cell_i_28 ( .A(A[28]), .B(B[28]), .p(P[28]), .g(G[28]) );
  PG_cell_3 PG_cell_i_29 ( .A(A[29]), .B(B[29]), .p(P[29]), .g(G[29]) );
  PG_cell_2 PG_cell_i_30 ( .A(A[30]), .B(B[30]), .p(P[30]), .g(G[30]) );
  PG_cell_1 PG_cell_i_31 ( .A(A[31]), .B(B[31]), .p(P[31]), .g(G[31]) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(tmp1) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_31 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_62 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_61 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_31 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_30 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_60 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_59 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_30 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_29 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_58 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_57 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_29 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_28 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_56 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_55 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_28 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_27 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_54 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_53 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_27 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_26 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_52 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_51 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_26 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_25 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_50 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_49 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_25 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_24 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_48 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_47 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_24 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_23 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_46 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_45 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_23 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_22 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_44 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_43 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_22 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_21 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_42 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_41 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_21 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_20 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_40 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_39 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_20 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_19 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_38 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_37 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_19 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_18 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_36 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_35 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_18 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_17 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_34 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_33 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_17 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_16 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_32 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_31 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_16 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_15 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_30 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_29 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_15 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_14 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_28 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_27 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_14 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_13 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_26 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_25 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_13 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_12 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_24 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_23 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_12 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_11 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_22 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_21 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_11 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_10 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_20 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_19 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_10 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_9 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_18 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_17 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_9 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_8 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_16 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_15 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_8 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_7 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_14 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_13 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_7 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_6 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_12 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_11 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_6 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_5 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_10 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_9 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_5 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_4 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_8 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_7 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_4 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_3 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_6 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_5 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_3 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_2 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_4 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_3 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_2 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_1 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n7, n8, n9;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n8) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n7), .A3(s_nq[0]), .ZN(n9) );
  t_ff_rst0_2 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_1 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_1 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n9), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n8), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n7) );
  NAND2_X1 U3 ( .A1(n9), .A2(n8), .ZN(s_toggle[1]) );
endmodule


module Mux_Bit_NBIT_Sel2_31 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_30 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_29 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_28 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_27 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_26 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_25 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_24 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_23 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_22 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_21 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_20 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_19 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_18 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_17 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_16 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_15 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_14 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_13 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_12 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_11 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_10 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_9 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_8 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_7 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_6 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_5 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_4 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_3 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_2 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module Mux_Bit_NBIT_Sel2_1 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n4, n6, n7, n8;

  OAI22_X1 U1 ( .A1(n8), .A2(n6), .B1(sel[1]), .B2(n7), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n8)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n7)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module D_FF_31 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_30 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_29 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_28 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_27 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_26 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_25 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_24 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_23 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_22 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_21 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_20 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_19 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_18 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_17 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_16 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_15 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_14 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_13 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_12 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_11 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_10 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_9 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_8 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_7 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_6 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_5 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_4 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_3 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_2 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module D_FF_1 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module ComparatorWithEnable_1055 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1054 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1053 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1052 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1051 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1050 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1049 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1048 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1047 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1046 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1045 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1044 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1043 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1042 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1041 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1040 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1039 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1038 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1037 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1036 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1035 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1034 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1033 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1032 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1031 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1030 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1029 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1028 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1027 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1026 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1025 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1024 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1023 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1022 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1021 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1020 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1019 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1018 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1017 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1016 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1015 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1014 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1013 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1012 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1011 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1010 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1009 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1008 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1007 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1006 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1005 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1004 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1003 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1002 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1001 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1000 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_999 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_998 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_997 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_996 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_995 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_994 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_993 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_992 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_991 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_990 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_989 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_988 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_987 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_986 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_985 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_984 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_983 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_982 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_981 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_980 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_979 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_978 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_977 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_976 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_975 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_974 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_973 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_972 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_971 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_970 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_969 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_968 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_967 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_966 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_965 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_964 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_963 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_962 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_961 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_960 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_959 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_958 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_957 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_956 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_955 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_954 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_953 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_952 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_951 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_950 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_949 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_948 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_947 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_946 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_945 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_944 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_943 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_942 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_941 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_940 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_939 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_938 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_937 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_936 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_935 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_934 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_933 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_932 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_931 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_930 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_929 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_928 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_927 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_926 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_925 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_924 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_923 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_922 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_921 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_920 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_919 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_918 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_917 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_916 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_915 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_914 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_913 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_912 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_911 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_910 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_909 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_908 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_907 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_906 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_905 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_904 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_903 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_902 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_901 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_900 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_899 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_898 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_897 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_896 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_895 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_894 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_893 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_892 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_891 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_890 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_889 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_888 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_887 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_886 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_885 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_884 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_883 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_882 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_881 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_880 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_879 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_878 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_877 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_876 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_875 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_874 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_873 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_872 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_871 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_870 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_869 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_868 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_867 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_866 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_865 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_864 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_863 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_862 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_861 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_860 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_859 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_858 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_857 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_856 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_855 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_854 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_853 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_852 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_851 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_850 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_849 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_848 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_847 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_846 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_845 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_844 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_843 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_842 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_841 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_840 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_839 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_838 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_837 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_836 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_835 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_834 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_833 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_832 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_831 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_830 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_829 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_828 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_827 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_826 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_825 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_824 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_823 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_822 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_821 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_820 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_819 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_818 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_817 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_816 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_815 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_814 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_813 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_812 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_811 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_810 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_809 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_808 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_807 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_806 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_805 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_804 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_803 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_802 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_801 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_800 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_799 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_798 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_797 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_796 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_795 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_794 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_793 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_792 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_791 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_790 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_789 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_788 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_787 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_786 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_785 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_784 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_783 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_782 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_781 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_780 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_779 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_778 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_777 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_776 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_775 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_774 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_773 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_772 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_771 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_770 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_769 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_768 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_767 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_766 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_765 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_764 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_763 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_762 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_761 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_760 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_759 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_758 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_757 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_756 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_755 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_754 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_753 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_752 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_751 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_750 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_749 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_748 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_747 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_746 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_745 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_744 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_743 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_742 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_741 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_740 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_739 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_738 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_737 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_736 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_735 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_734 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_733 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_732 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_731 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_730 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_729 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_728 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_727 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_726 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_725 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_724 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_723 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_722 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_721 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_720 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_719 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_718 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_717 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_716 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_715 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_714 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_713 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_712 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_711 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_710 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_709 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_708 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_707 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_706 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_705 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_704 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_703 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_702 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_701 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_700 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_699 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_698 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_697 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_696 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_695 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_694 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_693 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_692 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_691 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_690 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_689 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_688 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_687 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_686 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_685 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_684 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_683 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_682 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_681 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_680 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_679 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_678 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_677 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_676 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_675 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_674 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_673 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_672 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_671 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_670 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_669 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_668 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_667 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_666 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_665 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_664 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_663 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_662 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_661 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_660 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_659 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_658 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_657 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_656 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_655 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_654 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_653 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_652 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_651 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_650 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_649 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_648 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_647 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_646 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_645 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_644 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_643 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_642 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_641 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_640 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_639 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_638 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_637 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_636 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_635 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_634 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_633 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_632 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_631 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_630 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_629 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_628 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_627 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_626 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_625 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_624 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_623 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_622 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_621 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_620 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_619 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_618 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_617 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_616 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_615 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_614 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_613 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_612 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_611 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_610 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_609 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_608 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_607 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_606 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_605 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_604 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_603 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_602 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_601 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_600 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_599 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_598 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_597 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_596 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_595 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_594 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_593 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_592 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_591 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_590 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_589 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_588 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_587 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_586 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_585 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_584 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_583 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_582 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_581 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_580 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_579 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_578 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_577 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_576 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_575 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_574 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_573 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_572 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_571 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_570 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_569 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_568 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_567 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_566 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_565 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_564 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_563 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_562 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_561 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_560 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_559 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_558 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_557 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_556 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_555 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_554 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_553 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_552 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_551 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_550 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_549 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_548 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_547 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_546 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_545 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_544 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_543 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_542 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_541 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_540 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_539 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_538 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_537 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_536 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_535 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_534 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_533 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_532 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_531 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_530 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_529 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_528 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_527 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_526 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_525 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_524 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_523 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_522 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_521 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_520 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_519 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_518 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_517 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_516 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_515 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_514 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_513 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_512 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_511 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_510 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_509 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_508 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_507 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_506 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_505 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_504 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_503 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_502 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_501 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_500 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_499 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_498 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_497 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_496 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_495 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_494 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_493 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_492 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_491 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_490 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_489 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_488 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_487 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_486 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_485 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_484 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_483 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_482 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_481 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_480 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_479 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_478 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_477 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_476 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_475 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_474 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_473 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_472 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_471 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_470 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_469 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_468 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_467 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_466 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_465 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_464 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_463 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_462 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_461 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_460 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_459 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_458 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_457 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_456 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_455 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_454 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_453 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_452 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_451 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_450 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_449 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_448 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_447 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_446 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_445 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_444 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_443 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_442 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_441 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_440 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_439 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_438 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_437 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_436 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_435 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_434 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_433 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_432 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_431 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_430 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_429 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_428 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_427 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_426 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_425 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_424 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_423 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_422 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_421 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_420 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_419 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_418 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_417 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_416 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_415 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_414 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_413 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_412 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_411 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_410 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_409 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_408 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_407 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_406 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_405 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_404 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_403 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_402 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_401 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_400 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_399 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_398 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_397 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_396 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_395 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_394 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_393 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_392 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_391 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_390 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_389 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_388 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_387 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_386 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_385 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_384 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_383 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_382 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_381 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_380 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_379 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_378 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_377 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_376 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_375 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_374 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_373 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_372 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_371 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_370 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_369 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_368 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_367 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_366 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_365 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_364 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_363 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_362 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_361 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_360 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_359 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_358 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_357 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_356 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_355 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_354 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_353 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_352 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_351 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_350 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_349 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_348 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_347 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_346 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_345 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_344 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_343 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_342 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_341 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_340 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_339 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_338 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_337 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_336 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_335 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_334 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_333 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_332 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_331 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_330 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_329 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_328 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_327 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_326 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_325 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_324 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_323 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_322 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_321 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_320 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_319 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_318 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_317 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_316 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_315 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_314 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_313 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_312 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_311 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_310 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_309 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_308 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_307 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_306 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_305 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_304 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_303 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_302 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_301 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_300 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_299 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_298 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_297 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_296 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_295 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_294 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_293 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_292 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_291 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_290 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_289 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_288 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_287 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_286 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_285 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_284 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_283 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_282 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_281 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_280 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_279 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_278 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_277 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_276 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_275 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_274 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_273 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_272 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_271 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_270 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_269 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_268 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_267 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_266 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_265 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_264 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_263 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_262 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_261 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_260 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_259 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_258 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_257 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_256 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_255 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_254 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_253 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_252 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_251 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_250 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_249 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_248 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_247 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_246 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_245 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_244 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_243 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_242 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_241 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_240 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_239 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_238 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_237 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_236 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_235 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_234 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_233 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_232 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_231 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_230 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_229 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_228 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_227 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_226 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_225 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_224 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_223 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_222 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_221 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_220 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_219 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_218 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_217 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_216 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_215 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_214 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_213 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_212 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_211 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_210 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_209 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_208 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_207 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_206 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_205 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_204 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_203 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_202 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_201 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_200 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_199 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_198 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_197 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_196 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_195 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_194 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_193 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_192 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_191 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_190 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_189 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_188 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_187 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_186 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_185 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_184 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_183 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_182 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_181 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_180 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_179 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_178 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_177 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_176 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_175 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_174 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_173 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_172 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_171 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_170 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_169 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_168 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_167 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_166 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_165 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_164 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_163 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_162 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_161 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_160 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_159 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_158 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_157 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_156 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_155 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_154 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_153 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_152 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_151 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_150 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_149 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_148 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_147 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_146 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_145 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_144 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_143 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_142 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_141 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_140 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_139 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_138 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_137 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_136 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_135 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_134 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_133 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_132 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_131 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_130 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_129 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_128 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_127 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_126 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_125 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_124 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_123 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_122 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_121 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_120 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_119 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_118 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_117 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_116 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_115 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_114 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_113 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_112 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_111 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_110 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_109 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_108 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_107 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_106 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_105 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_104 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_103 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_102 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_101 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_100 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_99 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_98 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_97 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_96 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_95 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_94 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_93 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_92 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_91 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_90 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_89 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_88 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_87 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_86 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_85 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_84 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_83 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_82 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_81 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_80 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_79 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_78 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_77 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_76 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_75 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_74 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_73 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_72 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_71 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_70 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_69 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_68 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_67 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_66 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_65 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_64 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_63 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_62 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_61 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_60 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_59 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_58 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_57 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_56 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_55 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_54 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_53 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_52 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_51 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_50 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_49 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_48 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_47 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_46 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_45 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_44 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_43 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_42 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_41 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_40 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_39 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_38 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_37 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_36 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_35 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_34 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_33 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_32 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_31 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_30 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_29 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_28 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_27 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_26 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_25 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_24 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_23 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_22 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_21 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_20 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_19 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_18 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_17 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_16 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_15 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_14 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_13 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_12 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_11 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_10 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_9 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_8 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_7 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_6 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_5 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_4 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_3 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_2 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module ComparatorWithEnable_1 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n2;

  AND2_X1 U1 ( .A1(n2), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n2) );
endmodule


module CU_SatCounter_32 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_31 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_30 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_29 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_28 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_27 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_26 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_25 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_24 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_23 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_22 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_21 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_20 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_19 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_18 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_17 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_16 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_15 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_14 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_13 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_12 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_11 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_10 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_9 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_8 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_7 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_6 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_5 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_4 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_3 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_2 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module CU_SatCounter_1 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n8, n10, n11, n12, n13, n14;
  assign UDC_clk = CU_clk;

  INV_X1 U3 ( .A(n14), .ZN(UDC_reset) );
  AOI21_X1 U4 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n14) );
  NOR3_X1 U5 ( .A1(CU_TcMax), .A2(n12), .A3(n8), .ZN(UDC_Ud) );
  OR2_X1 U6 ( .A1(n13), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U7 ( .A1(n12), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n13) );
  NAND4_X1 U8 ( .A1(CU_update), .A2(CU_enable), .A3(n11), .A4(n10), .ZN(n12)
         );
  INV_X1 U9 ( .A(CU_loadDefault), .ZN(n11) );
  INV_X1 U10 ( .A(CU_Ud), .ZN(n8) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module Enable_Interface_NBIT_DATA32_3 ( EI_datain, EI_enable, EI_dataout );
  input [31:0] EI_datain;
  output [31:0] EI_dataout;
  input EI_enable;
  wire   n1, n2, n3;

  AND2_X1 U1 ( .A1(EI_datain[31]), .A2(n3), .ZN(EI_dataout[31]) );
  AND2_X1 U2 ( .A1(EI_datain[26]), .A2(n2), .ZN(EI_dataout[26]) );
  AND2_X1 U3 ( .A1(EI_datain[30]), .A2(n2), .ZN(EI_dataout[30]) );
  AND2_X1 U4 ( .A1(EI_datain[27]), .A2(n2), .ZN(EI_dataout[27]) );
  AND2_X1 U5 ( .A1(EI_datain[21]), .A2(n2), .ZN(EI_dataout[21]) );
  AND2_X1 U6 ( .A1(EI_datain[24]), .A2(n2), .ZN(EI_dataout[24]) );
  AND2_X1 U7 ( .A1(EI_datain[18]), .A2(n1), .ZN(EI_dataout[18]) );
  AND2_X1 U8 ( .A1(EI_datain[15]), .A2(n1), .ZN(EI_dataout[15]) );
  AND2_X1 U9 ( .A1(EI_datain[28]), .A2(n2), .ZN(EI_dataout[28]) );
  AND2_X1 U10 ( .A1(EI_datain[22]), .A2(n2), .ZN(EI_dataout[22]) );
  AND2_X1 U11 ( .A1(EI_datain[20]), .A2(n2), .ZN(EI_dataout[20]) );
  AND2_X1 U12 ( .A1(EI_datain[17]), .A2(n1), .ZN(EI_dataout[17]) );
  AND2_X1 U13 ( .A1(EI_datain[29]), .A2(n2), .ZN(EI_dataout[29]) );
  AND2_X1 U14 ( .A1(EI_datain[23]), .A2(n2), .ZN(EI_dataout[23]) );
  AND2_X1 U15 ( .A1(EI_datain[16]), .A2(n1), .ZN(EI_dataout[16]) );
  AND2_X1 U16 ( .A1(EI_datain[19]), .A2(n1), .ZN(EI_dataout[19]) );
  AND2_X1 U17 ( .A1(EI_datain[25]), .A2(n2), .ZN(EI_dataout[25]) );
  AND2_X1 U18 ( .A1(EI_datain[12]), .A2(n1), .ZN(EI_dataout[12]) );
  AND2_X1 U19 ( .A1(n3), .A2(EI_datain[9]), .ZN(EI_dataout[9]) );
  AND2_X1 U20 ( .A1(EI_datain[6]), .A2(n3), .ZN(EI_dataout[6]) );
  AND2_X1 U21 ( .A1(EI_datain[10]), .A2(n1), .ZN(EI_dataout[10]) );
  AND2_X1 U22 ( .A1(EI_datain[13]), .A2(n1), .ZN(EI_dataout[13]) );
  AND2_X1 U23 ( .A1(EI_datain[11]), .A2(n1), .ZN(EI_dataout[11]) );
  AND2_X1 U24 ( .A1(EI_datain[14]), .A2(n1), .ZN(EI_dataout[14]) );
  AND2_X1 U25 ( .A1(EI_datain[8]), .A2(n3), .ZN(EI_dataout[8]) );
  AND2_X1 U26 ( .A1(EI_datain[7]), .A2(n3), .ZN(EI_dataout[7]) );
  AND2_X1 U27 ( .A1(EI_datain[1]), .A2(n1), .ZN(EI_dataout[1]) );
  AND2_X1 U28 ( .A1(EI_datain[3]), .A2(n3), .ZN(EI_dataout[3]) );
  AND2_X1 U29 ( .A1(EI_datain[0]), .A2(n1), .ZN(EI_dataout[0]) );
  AND2_X1 U30 ( .A1(EI_datain[2]), .A2(n2), .ZN(EI_dataout[2]) );
  AND2_X1 U31 ( .A1(EI_datain[4]), .A2(n3), .ZN(EI_dataout[4]) );
  AND2_X1 U32 ( .A1(EI_datain[5]), .A2(n3), .ZN(EI_dataout[5]) );
  CLKBUF_X1 U33 ( .A(EI_enable), .Z(n2) );
  CLKBUF_X1 U34 ( .A(EI_enable), .Z(n3) );
  CLKBUF_X1 U35 ( .A(EI_enable), .Z(n1) );
endmodule


module Enable_Interface_NBIT_DATA32_2 ( EI_datain, EI_enable, EI_dataout );
  input [31:0] EI_datain;
  output [31:0] EI_dataout;
  input EI_enable;
  wire   net142017, net142015, net142013;

  AND2_X2 U1 ( .A1(EI_datain[0]), .A2(net142013), .ZN(EI_dataout[0]) );
  BUF_X2 U2 ( .A(EI_enable), .Z(net142013) );
  CLKBUF_X1 U3 ( .A(EI_enable), .Z(net142015) );
  CLKBUF_X1 U4 ( .A(EI_enable), .Z(net142017) );
  AND2_X2 U5 ( .A1(EI_datain[1]), .A2(net142013), .ZN(EI_dataout[1]) );
  AND2_X2 U6 ( .A1(EI_datain[2]), .A2(net142015), .ZN(EI_dataout[2]) );
  AND2_X1 U7 ( .A1(EI_datain[3]), .A2(net142017), .ZN(EI_dataout[3]) );
  AND2_X1 U8 ( .A1(EI_datain[4]), .A2(net142017), .ZN(EI_dataout[4]) );
  AND2_X1 U9 ( .A1(EI_datain[5]), .A2(net142017), .ZN(EI_dataout[5]) );
  AND2_X1 U10 ( .A1(EI_datain[6]), .A2(net142017), .ZN(EI_dataout[6]) );
  AND2_X1 U11 ( .A1(EI_datain[10]), .A2(net142013), .ZN(EI_dataout[10]) );
  AND2_X1 U12 ( .A1(EI_datain[11]), .A2(net142013), .ZN(EI_dataout[11]) );
  AND2_X1 U13 ( .A1(EI_datain[12]), .A2(net142013), .ZN(EI_dataout[12]) );
  AND2_X1 U14 ( .A1(EI_datain[15]), .A2(net142013), .ZN(EI_dataout[15]) );
  AND2_X1 U15 ( .A1(EI_datain[13]), .A2(net142013), .ZN(EI_dataout[13]) );
  AND2_X1 U16 ( .A1(EI_datain[16]), .A2(net142013), .ZN(EI_dataout[16]) );
  AND2_X1 U17 ( .A1(EI_datain[14]), .A2(net142013), .ZN(EI_dataout[14]) );
  AND2_X1 U18 ( .A1(EI_datain[17]), .A2(net142013), .ZN(EI_dataout[17]) );
  AND2_X1 U19 ( .A1(EI_datain[18]), .A2(net142013), .ZN(EI_dataout[18]) );
  AND2_X1 U20 ( .A1(EI_datain[19]), .A2(net142013), .ZN(EI_dataout[19]) );
  AND2_X1 U21 ( .A1(EI_datain[20]), .A2(net142015), .ZN(EI_dataout[20]) );
  AND2_X1 U22 ( .A1(EI_datain[21]), .A2(net142015), .ZN(EI_dataout[21]) );
  AND2_X1 U23 ( .A1(EI_datain[22]), .A2(net142015), .ZN(EI_dataout[22]) );
  AND2_X1 U24 ( .A1(net142017), .A2(EI_datain[9]), .ZN(EI_dataout[9]) );
  AND2_X1 U25 ( .A1(EI_datain[7]), .A2(net142017), .ZN(EI_dataout[7]) );
  AND2_X1 U26 ( .A1(EI_datain[8]), .A2(net142017), .ZN(EI_dataout[8]) );
  AND2_X1 U27 ( .A1(EI_datain[23]), .A2(net142015), .ZN(EI_dataout[23]) );
  AND2_X1 U28 ( .A1(EI_datain[24]), .A2(net142015), .ZN(EI_dataout[24]) );
  AND2_X1 U29 ( .A1(EI_datain[25]), .A2(net142015), .ZN(EI_dataout[25]) );
  AND2_X1 U30 ( .A1(EI_datain[26]), .A2(net142015), .ZN(EI_dataout[26]) );
  AND2_X1 U31 ( .A1(EI_datain[27]), .A2(net142015), .ZN(EI_dataout[27]) );
  AND2_X1 U32 ( .A1(EI_datain[28]), .A2(net142015), .ZN(EI_dataout[28]) );
  AND2_X1 U33 ( .A1(EI_datain[29]), .A2(net142015), .ZN(EI_dataout[29]) );
  AND2_X1 U34 ( .A1(EI_datain[30]), .A2(net142015), .ZN(EI_dataout[30]) );
  AND2_X1 U35 ( .A1(EI_datain[31]), .A2(net142017), .ZN(EI_dataout[31]) );
endmodule


module Enable_Interface_NBIT_DATA32_1 ( EI_datain, EI_enable, EI_dataout );
  input [31:0] EI_datain;
  output [31:0] EI_dataout;
  input EI_enable;
  wire   n1, n2, n3;

  AND2_X2 U8 ( .A1(EI_datain[31]), .A2(n3), .ZN(EI_dataout[31]) );
  AND2_X2 U18 ( .A1(EI_datain[22]), .A2(n2), .ZN(EI_dataout[22]) );
  AND2_X2 U1 ( .A1(EI_datain[29]), .A2(n2), .ZN(EI_dataout[29]) );
  AND2_X1 U2 ( .A1(EI_datain[1]), .A2(n1), .ZN(EI_dataout[1]) );
  AND2_X1 U3 ( .A1(EI_datain[2]), .A2(n2), .ZN(EI_dataout[2]) );
  AND2_X1 U4 ( .A1(EI_datain[3]), .A2(n3), .ZN(EI_dataout[3]) );
  AND2_X1 U5 ( .A1(EI_datain[4]), .A2(n3), .ZN(EI_dataout[4]) );
  AND2_X1 U6 ( .A1(EI_datain[5]), .A2(n3), .ZN(EI_dataout[5]) );
  AND2_X1 U7 ( .A1(EI_datain[6]), .A2(n3), .ZN(EI_dataout[6]) );
  AND2_X1 U9 ( .A1(EI_datain[7]), .A2(n3), .ZN(EI_dataout[7]) );
  AND2_X1 U10 ( .A1(EI_datain[8]), .A2(n3), .ZN(EI_dataout[8]) );
  AND2_X1 U11 ( .A1(n3), .A2(EI_datain[9]), .ZN(EI_dataout[9]) );
  AND2_X1 U12 ( .A1(EI_datain[10]), .A2(n1), .ZN(EI_dataout[10]) );
  AND2_X1 U13 ( .A1(EI_datain[11]), .A2(n1), .ZN(EI_dataout[11]) );
  AND2_X1 U14 ( .A1(EI_datain[12]), .A2(n1), .ZN(EI_dataout[12]) );
  AND2_X1 U15 ( .A1(EI_datain[13]), .A2(n1), .ZN(EI_dataout[13]) );
  AND2_X1 U16 ( .A1(EI_datain[14]), .A2(n1), .ZN(EI_dataout[14]) );
  AND2_X1 U17 ( .A1(EI_datain[15]), .A2(n1), .ZN(EI_dataout[15]) );
  AND2_X1 U19 ( .A1(EI_datain[16]), .A2(n1), .ZN(EI_dataout[16]) );
  AND2_X1 U20 ( .A1(EI_datain[17]), .A2(n1), .ZN(EI_dataout[17]) );
  AND2_X1 U21 ( .A1(EI_datain[18]), .A2(n1), .ZN(EI_dataout[18]) );
  AND2_X1 U22 ( .A1(EI_datain[19]), .A2(n1), .ZN(EI_dataout[19]) );
  AND2_X1 U23 ( .A1(EI_datain[20]), .A2(n2), .ZN(EI_dataout[20]) );
  AND2_X1 U24 ( .A1(EI_datain[21]), .A2(n2), .ZN(EI_dataout[21]) );
  AND2_X1 U25 ( .A1(EI_datain[23]), .A2(n2), .ZN(EI_dataout[23]) );
  AND2_X1 U26 ( .A1(EI_datain[24]), .A2(n2), .ZN(EI_dataout[24]) );
  AND2_X2 U27 ( .A1(EI_datain[25]), .A2(n2), .ZN(EI_dataout[25]) );
  AND2_X2 U28 ( .A1(EI_datain[26]), .A2(n2), .ZN(EI_dataout[26]) );
  AND2_X2 U29 ( .A1(EI_datain[27]), .A2(n2), .ZN(EI_dataout[27]) );
  AND2_X2 U30 ( .A1(EI_datain[30]), .A2(n2), .ZN(EI_dataout[30]) );
  AND2_X2 U31 ( .A1(EI_datain[28]), .A2(n2), .ZN(EI_dataout[28]) );
  CLKBUF_X1 U32 ( .A(EI_enable), .Z(n1) );
  CLKBUF_X3 U33 ( .A(EI_enable), .Z(n2) );
  AND2_X1 U34 ( .A1(EI_datain[0]), .A2(n1), .ZN(EI_dataout[0]) );
  CLKBUF_X3 U35 ( .A(EI_enable), .Z(n3) );
endmodule


module NRegister_N5_2 ( clk, reset, data_in, enable, load, data_out );
  input [4:0] data_in;
  output [4:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, net110627, net110628, net110629, net110630,
         net110631, n8, n9, n10, n11, n12, n13, n16, n17;

  DFFR_X1 \data_out_reg[4]  ( .D(n2), .CK(clk), .RN(n8), .Q(data_out[4]), .QN(
        net110631) );
  DFFR_X1 \data_out_reg[3]  ( .D(n4), .CK(clk), .RN(n8), .Q(data_out[3]), .QN(
        net110630) );
  DFFR_X1 \data_out_reg[2]  ( .D(n5), .CK(clk), .RN(n8), .Q(data_out[2]), .QN(
        net110629) );
  DFFR_X1 \data_out_reg[1]  ( .D(n6), .CK(clk), .RN(n8), .Q(data_out[1]), .QN(
        net110628) );
  DFFR_X1 \data_out_reg[0]  ( .D(n7), .CK(clk), .RN(n8), .Q(data_out[0]), .QN(
        net110627) );
  INV_X1 U3 ( .A(n17), .ZN(n13) );
  NAND2_X1 U4 ( .A1(load), .A2(enable), .ZN(n17) );
  OAI22_X1 U5 ( .A1(n17), .A2(n16), .B1(net110627), .B2(n13), .ZN(n7) );
  INV_X1 U6 ( .A(data_in[0]), .ZN(n16) );
  OAI22_X1 U7 ( .A1(n17), .A2(n12), .B1(net110628), .B2(n13), .ZN(n6) );
  INV_X1 U8 ( .A(data_in[1]), .ZN(n12) );
  OAI22_X1 U9 ( .A1(n17), .A2(n11), .B1(net110629), .B2(n13), .ZN(n5) );
  INV_X1 U10 ( .A(data_in[2]), .ZN(n11) );
  OAI22_X1 U11 ( .A1(n17), .A2(n10), .B1(net110630), .B2(n13), .ZN(n4) );
  INV_X1 U12 ( .A(data_in[3]), .ZN(n10) );
  OAI22_X1 U13 ( .A1(n17), .A2(n9), .B1(net110631), .B2(n13), .ZN(n2) );
  INV_X1 U14 ( .A(data_in[4]), .ZN(n9) );
  INV_X1 U15 ( .A(reset), .ZN(n8) );
endmodule


module NRegister_N5_1 ( clk, reset, data_in, enable, load, data_out );
  input [4:0] data_in;
  output [4:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n3, n4, n5, n6, n7, net110627, net110628, net110629, net110630,
         net110631, n8, n9, n10, n11, n12, n13, n15;

  DFFR_X1 \data_out_reg[4]  ( .D(n2), .CK(clk), .RN(n3), .Q(data_out[4]), .QN(
        net110631) );
  DFFR_X1 \data_out_reg[3]  ( .D(n4), .CK(clk), .RN(n3), .Q(data_out[3]), .QN(
        net110630) );
  DFFR_X1 \data_out_reg[2]  ( .D(n5), .CK(clk), .RN(n3), .Q(data_out[2]), .QN(
        net110629) );
  DFFR_X1 \data_out_reg[0]  ( .D(n7), .CK(clk), .RN(n3), .Q(data_out[0]), .QN(
        net110627) );
  DFFR_X2 \data_out_reg[1]  ( .D(n6), .CK(clk), .RN(n3), .Q(data_out[1]), .QN(
        net110628) );
  INV_X1 U3 ( .A(n15), .ZN(n12) );
  OAI22_X1 U4 ( .A1(n15), .A2(n13), .B1(net110627), .B2(n12), .ZN(n7) );
  INV_X1 U5 ( .A(data_in[0]), .ZN(n13) );
  OAI22_X1 U6 ( .A1(n15), .A2(n9), .B1(net110630), .B2(n12), .ZN(n4) );
  INV_X1 U7 ( .A(data_in[3]), .ZN(n9) );
  OAI22_X1 U8 ( .A1(n15), .A2(n10), .B1(net110629), .B2(n12), .ZN(n5) );
  INV_X1 U9 ( .A(data_in[2]), .ZN(n10) );
  OAI22_X1 U10 ( .A1(n15), .A2(n8), .B1(net110631), .B2(n12), .ZN(n2) );
  INV_X1 U11 ( .A(data_in[4]), .ZN(n8) );
  NAND2_X1 U12 ( .A1(load), .A2(enable), .ZN(n15) );
  INV_X1 U13 ( .A(reset), .ZN(n3) );
  OAI22_X1 U14 ( .A1(n11), .A2(n15), .B1(net110628), .B2(n12), .ZN(n6) );
  INV_X1 U15 ( .A(data_in[1]), .ZN(n11) );
endmodule


module PropagateCarryLookahead_N32_1 ( A, B, Cin, Sum, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Sum;
  input Cin;
  output Cout;

  wire   [31:0] s_G1;
  wire   [31:0] s_P1;
  wire   [31:0] s_G2;
  wire   [31:0] s_P2;
  wire   SYNOPSYS_UNCONNECTED__0;

  PG_network_N32_2 PG ( .A(A), .B(B), .c_in(1'b0), .G(s_G1), .P({s_P1[31:1], 
        SYNOPSYS_UNCONNECTED__0}) );
  Carry_Network_N32_1 CN ( .G(s_G1), .P({s_P1[31:1], 1'b0}), .Cin(Cin), .Cout(
        Cout), .Gout(s_G2), .Pout(s_P2) );
  Sum_Network_N32_1 SN ( .G(s_G2), .P(s_P2), .S(Sum) );
endmodule


module SAT_Counter_BTB_N3_31 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_31 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_31 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_30 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_30 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_30 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_29 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_29 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_29 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_28 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_28 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_28 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_27 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_27 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_27 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_26 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_26 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_26 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_25 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_25 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_25 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_24 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_24 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_24 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_23 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_23 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_23 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_22 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_22 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_22 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_21 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_21 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_21 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_20 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_20 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_20 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_19 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_19 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_19 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_18 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_18 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_18 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_17 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_17 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_17 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_16 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_16 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_16 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_15 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_15 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_15 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_14 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_14 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_14 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_13 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_13 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_13 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_12 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_12 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_12 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_11 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_11 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_11 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_10 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_10 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), 
        .UDC_CLK(s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_10 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_9 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_9 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), .UDC_CLK(
        s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_9 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_8 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_8 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), .UDC_CLK(
        s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_8 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_7 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_7 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), .UDC_CLK(
        s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_7 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_6 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_6 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), .UDC_CLK(
        s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_6 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_5 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_5 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), .UDC_CLK(
        s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_5 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_4 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_4 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), .UDC_CLK(
        s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_4 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_3 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_3 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), .UDC_CLK(
        s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_3 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_2 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_2 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), .UDC_CLK(
        s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_2 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module SAT_Counter_BTB_N3_1 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_1 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), .UDC_CLK(
        s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_1 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module ORGate_NX1_N32_1 ( A, B, Y );
  input [31:0] A;
  input [31:0] B;
  output Y;
  wire   n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34,
         n35, n36, n37, n38, n39, n40, n41, n42;

  AND2_X1 U1 ( .A1(n33), .A2(n31), .ZN(n21) );
  NAND4_X1 U2 ( .A1(n22), .A2(n23), .A3(n24), .A4(n25), .ZN(Y) );
  AND3_X1 U3 ( .A1(n34), .A2(n32), .A3(n21), .ZN(n22) );
  AND4_X1 U4 ( .A1(n30), .A2(n29), .A3(n28), .A4(n27), .ZN(n23) );
  AND4_X1 U5 ( .A1(n38), .A2(n37), .A3(n36), .A4(n35), .ZN(n24) );
  AND4_X1 U6 ( .A1(n42), .A2(n41), .A3(n40), .A4(n39), .ZN(n25) );
  NOR4_X1 U7 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n32) );
  NOR4_X1 U8 ( .A1(A[30]), .A2(A[2]), .A3(A[29]), .A4(A[28]), .ZN(n29) );
  OR3_X1 U9 ( .A1(A[10]), .A2(A[11]), .A3(A[12]), .ZN(n26) );
  NOR4_X1 U10 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n27) );
  NOR4_X1 U11 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n30) );
  NOR4_X1 U12 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n28) );
  NOR4_X1 U13 ( .A1(B[9]), .A2(B[8]), .A3(B[7]), .A4(B[6]), .ZN(n35) );
  NOR4_X1 U14 ( .A1(B[23]), .A2(B[22]), .A3(B[21]), .A4(B[20]), .ZN(n39) );
  NOR4_X1 U15 ( .A1(B[5]), .A2(B[4]), .A3(B[3]), .A4(B[31]), .ZN(n36) );
  NOR4_X1 U16 ( .A1(B[1]), .A2(B[19]), .A3(B[18]), .A4(B[17]), .ZN(n40) );
  NOR4_X1 U17 ( .A1(B[30]), .A2(B[2]), .A3(B[29]), .A4(B[28]), .ZN(n37) );
  NOR4_X1 U18 ( .A1(B[16]), .A2(B[15]), .A3(B[14]), .A4(B[13]), .ZN(n41) );
  NOR4_X1 U19 ( .A1(B[27]), .A2(B[26]), .A3(B[25]), .A4(B[24]), .ZN(n38) );
  NOR4_X1 U20 ( .A1(B[12]), .A2(B[11]), .A3(B[10]), .A4(B[0]), .ZN(n42) );
  NOR2_X1 U21 ( .A1(A[0]), .A2(n26), .ZN(n34) );
  NOR4_X1 U22 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n31) );
  NOR4_X1 U23 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n33) );
endmodule


module NComparatorWithEnable_NBIT32_32 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_1024 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_1023 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_1022 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_1021 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_1020 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_1019 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_1018 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_1017 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_1016 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_1015 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_1014 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_1013 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_1012 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_1011 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_1010 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_1009 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_1008 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_1007 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_1006 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_1005 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_1004 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_1003 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_1002 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_1001 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_1000 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_999 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_998 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_997 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_996 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_995 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_994 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_993 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_31 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_992 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_991 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_990 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_989 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_988 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_987 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_986 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_985 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_984 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_983 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_982 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_981 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_980 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_979 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_978 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_977 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_976 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_975 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_974 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_973 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_972 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_971 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_970 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_969 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_968 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_967 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_966 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_965 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_964 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_963 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_962 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_961 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_30 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_960 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_959 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_958 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_957 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_956 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_955 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_954 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_953 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_952 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_951 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_950 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_949 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_948 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_947 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_946 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_945 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_944 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_943 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_942 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_941 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_940 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_939 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_938 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_937 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_936 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_935 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_934 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_933 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_932 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_931 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_930 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_929 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_29 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_928 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_927 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_926 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_925 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_924 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_923 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_922 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_921 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_920 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_919 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_918 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_917 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_916 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_915 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_914 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_913 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_912 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_911 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_910 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_909 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_908 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_907 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_906 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_905 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_904 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_903 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_902 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_901 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_900 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_899 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_898 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_897 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_28 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_896 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_895 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_894 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_893 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_892 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_891 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_890 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_889 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_888 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_887 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_886 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_885 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_884 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_883 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_882 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_881 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_880 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_879 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_878 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_877 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_876 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_875 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_874 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_873 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_872 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_871 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_870 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_869 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_868 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_867 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_866 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_865 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_27 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_864 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_863 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_862 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_861 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_860 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_859 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_858 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_857 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_856 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_855 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_854 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_853 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_852 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_851 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_850 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_849 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_848 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_847 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_846 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_845 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_844 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_843 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_842 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_841 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_840 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_839 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_838 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_837 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_836 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_835 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_834 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_833 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_26 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_832 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_831 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_830 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_829 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_828 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_827 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_826 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_825 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_824 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_823 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_822 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_821 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_820 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_819 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_818 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_817 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_816 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_815 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_814 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_813 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_812 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_811 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_810 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_809 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_808 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_807 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_806 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_805 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_804 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_803 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_802 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_801 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_25 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_800 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_799 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_798 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_797 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_796 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_795 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_794 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_793 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_792 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_791 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_790 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_789 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_788 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_787 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_786 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_785 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_784 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_783 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_782 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_781 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_780 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_779 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_778 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_777 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_776 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_775 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_774 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_773 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_772 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_771 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_770 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_769 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_24 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_768 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_767 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_766 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_765 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_764 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_763 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_762 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_761 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_760 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_759 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_758 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_757 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_756 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_755 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_754 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_753 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_752 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_751 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_750 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_749 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_748 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_747 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_746 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_745 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_744 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_743 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_742 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_741 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_740 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_739 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_738 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_737 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_23 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_736 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_735 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_734 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_733 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_732 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_731 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_730 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_729 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_728 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_727 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_726 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_725 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_724 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_723 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_722 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_721 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_720 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_719 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_718 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_717 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_716 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_715 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_714 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_713 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_712 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_711 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_710 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_709 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_708 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_707 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_706 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_705 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_22 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_704 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_703 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_702 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_701 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_700 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_699 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_698 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_697 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_696 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_695 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_694 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_693 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_692 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_691 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_690 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_689 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_688 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_687 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_686 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_685 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_684 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_683 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_682 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_681 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_680 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_679 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_678 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_677 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_676 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_675 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_674 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_673 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_21 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_672 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_671 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_670 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_669 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_668 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_667 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_666 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_665 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_664 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_663 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_662 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_661 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_660 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_659 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_658 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_657 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_656 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_655 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_654 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_653 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_652 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_651 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_650 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_649 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_648 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_647 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_646 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_645 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_644 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_643 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_642 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_641 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_20 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_640 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_639 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_638 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_637 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_636 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_635 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_634 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_633 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_632 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_631 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_630 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_629 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_628 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_627 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_626 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_625 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_624 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_623 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_622 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_621 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_620 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_619 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_618 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_617 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_616 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_615 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_614 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_613 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_612 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_611 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_610 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_609 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_19 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_608 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_607 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_606 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_605 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_604 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_603 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_602 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_601 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_600 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_599 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_598 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_597 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_596 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_595 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_594 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_593 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_592 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_591 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_590 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_589 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_588 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_587 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_586 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_585 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_584 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_583 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_582 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_581 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_580 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_579 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_578 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_577 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_18 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_576 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_575 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_574 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_573 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_572 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_571 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_570 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_569 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_568 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_567 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_566 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_565 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_564 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_563 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_562 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_561 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_560 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_559 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_558 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_557 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_556 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_555 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_554 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_553 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_552 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_551 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_550 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_549 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_548 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_547 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_546 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_545 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_17 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_544 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_543 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_542 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_541 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_540 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_539 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_538 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_537 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_536 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_535 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_534 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_533 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_532 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_531 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_530 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_529 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_528 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_527 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_526 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_525 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_524 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_523 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_522 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_521 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_520 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_519 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_518 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_517 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_516 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_515 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_514 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_513 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_16 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_512 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_511 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_510 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_509 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_508 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_507 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_506 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_505 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_504 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_503 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_502 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_501 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_500 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_499 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_498 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_497 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_496 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_495 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_494 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_493 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_492 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_491 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_490 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_489 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_488 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_487 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_486 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_485 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_484 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_483 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_482 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_481 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_15 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_480 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_479 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_478 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_477 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_476 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_475 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_474 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_473 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_472 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_471 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_470 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_469 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_468 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_467 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_466 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_465 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_464 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_463 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_462 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_461 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_460 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_459 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_458 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_457 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_456 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_455 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_454 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_453 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_452 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_451 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_450 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_449 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_14 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_448 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_447 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_446 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_445 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_444 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_443 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_442 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_441 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_440 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_439 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_438 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_437 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_436 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_435 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_434 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_433 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_432 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_431 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_430 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_429 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_428 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_427 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_426 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_425 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_424 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_423 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_422 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_421 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_420 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_419 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_418 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_417 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_13 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_416 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_415 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_414 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_413 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_412 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_411 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_410 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_409 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_408 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_407 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_406 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_405 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_404 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_403 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_402 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_401 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_400 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_399 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_398 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_397 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_396 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_395 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_394 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_393 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_392 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_391 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_390 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_389 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_388 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_387 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_386 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_385 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_12 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_384 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_383 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_382 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_381 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_380 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_379 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_378 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_377 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_376 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_375 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_374 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_373 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_372 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_371 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_370 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_369 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_368 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_367 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_366 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_365 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_364 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_363 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_362 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_361 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_360 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_359 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_358 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_357 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_356 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_355 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_354 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_353 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_11 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_352 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_351 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_350 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_349 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_348 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_347 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_346 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_345 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_344 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_343 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_342 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_341 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_340 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_339 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_338 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_337 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_336 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_335 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_334 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_333 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_332 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_331 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_330 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_329 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_328 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_327 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_326 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_325 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_324 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_323 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_322 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_321 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_10 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_320 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_319 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_318 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_317 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_316 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_315 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_314 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_313 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_312 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_311 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_310 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_309 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_308 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_307 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_306 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_305 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_304 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_303 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_302 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_301 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_300 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_299 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_298 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_297 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_296 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_295 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_294 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_293 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_292 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_291 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_290 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_289 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_9 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_288 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_287 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_286 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_285 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_284 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_283 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_282 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_281 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_280 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_279 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_278 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_277 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_276 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_275 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_274 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_273 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_272 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_271 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_270 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_269 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_268 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_267 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_266 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_265 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_264 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_263 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_262 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_261 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_260 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_259 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_258 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_257 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_8 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_256 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_255 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_254 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_253 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_252 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_251 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_250 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_249 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_248 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_247 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_246 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_245 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_244 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_243 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_242 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_241 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_240 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_239 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_238 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_237 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_236 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_235 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_234 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_233 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_232 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_231 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_230 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_229 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_228 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_227 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_226 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_225 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_7 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_224 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_223 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_222 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_221 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_220 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_219 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_218 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_217 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_216 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_215 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_214 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_213 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_212 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_211 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_210 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_209 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_208 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_207 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_206 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_205 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_204 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_203 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_202 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_201 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_200 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_199 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_198 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_197 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_196 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_195 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_194 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_193 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_6 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_192 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_191 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_190 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_189 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_188 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_187 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_186 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_185 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_184 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_183 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_182 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_181 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_180 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_179 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_178 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_177 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_176 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_175 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_174 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_173 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_172 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_171 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_170 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_169 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_168 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_167 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_166 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_165 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_164 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_163 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_162 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_161 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_5 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_160 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_159 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_158 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_157 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_156 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_155 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_154 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_153 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_152 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_151 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_150 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_149 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_148 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_147 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_146 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_145 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_144 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_143 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_142 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_141 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_140 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_139 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_138 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_137 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_136 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_135 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_134 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_133 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_132 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_131 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_130 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_129 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_4 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_128 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_127 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_126 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_125 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_124 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_123 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_122 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_121 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_120 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_119 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_118 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_117 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_116 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_115 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_114 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_113 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_112 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_111 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_110 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_109 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_108 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_107 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_106 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_105 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_104 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_103 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_102 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_101 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_100 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_99 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_98 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_97 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_3 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_96 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_95 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_94 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_93 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_92 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_91 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_90 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_89 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_88 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_87 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_86 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_85 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_84 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_83 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_82 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_81 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_80 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_79 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_78 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_77 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_76 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_75 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_74 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_73 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_72 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_71 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_70 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_69 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_68 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_67 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_66 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_65 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module NComparatorWithEnable_NBIT32_2 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;
  assign n3 = Enable;

  ComparatorWithEnable_64 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n14), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_63 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_62 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_61 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_60 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_59 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_58 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_57 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_56 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_55 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_54 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_53 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_52 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n15), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_51 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_50 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_49 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_48 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_47 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_46 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_45 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_44 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_43 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_42 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_41 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_40 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n16), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_39 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_38 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_37 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_36 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_35 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_34 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_33 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  AND2_X1 U4 ( .A1(n26), .A2(n25), .ZN(ComparatorBit) );
  NOR4_X1 U5 ( .A1(n20), .A2(n19), .A3(n18), .A4(n17), .ZN(n26) );
  NOR4_X1 U6 ( .A1(n24), .A2(n23), .A3(n22), .A4(n21), .ZN(n25) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n20) );
  NAND4_X1 U8 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n21) );
  NAND4_X1 U9 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n17) );
  NAND4_X1 U10 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(
        \matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n22) );
  NAND4_X1 U11 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n18) );
  NAND4_X1 U12 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n23) );
  NAND4_X1 U13 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n19) );
  NAND4_X1 U14 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n24) );
endmodule


module Mux_1Bit_2X1_7 ( port0, port1, sel, portY );
  input port0, port1, sel;
  output portY;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(portY) );
  AOI22_X1 U2 ( .A1(port0), .A2(n1), .B1(sel), .B2(port1), .ZN(n2) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module Mux_1Bit_2X1_5 ( port0, port1, sel, portY );
  input port0, port1, sel;
  output portY;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(portY) );
  AOI22_X1 U2 ( .A1(port0), .A2(n1), .B1(sel), .B2(port1), .ZN(n2) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module Mux_1Bit_2X1_3 ( port0, port1, sel, portY );
  input port0, port1, sel;
  output portY;
  wire   n1, n2, n3;

  NAND2_X1 U1 ( .A1(port0), .A2(n1), .ZN(n2) );
  NAND2_X1 U2 ( .A1(port1), .A2(sel), .ZN(n3) );
  NAND2_X1 U3 ( .A1(n2), .A2(n3), .ZN(portY) );
  INV_X1 U4 ( .A(sel), .ZN(n1) );
endmodule


module Mux_1Bit_2X1_2 ( port0, port1, sel, portY );
  input port0, port1, sel;
  output portY;
  wire   n1, n2, n5;

  NAND2_X1 U1 ( .A1(port0), .A2(n5), .ZN(n1) );
  NAND2_X1 U2 ( .A1(port1), .A2(sel), .ZN(n2) );
  NAND2_X1 U3 ( .A1(n2), .A2(n1), .ZN(portY) );
  INV_X1 U4 ( .A(sel), .ZN(n5) );
endmodule


module Mux_1Bit_2X1_1 ( port0, port1, sel, portY );
  input port0, port1, sel;
  output portY;
  wire   n1, n2;

  INV_X1 U1 ( .A(n2), .ZN(portY) );
  INV_X1 U2 ( .A(sel), .ZN(n1) );
  AOI22_X1 U3 ( .A1(port0), .A2(n1), .B1(port1), .B2(sel), .ZN(n2) );
endmodule


module Mux_NBit_2x1_NBIT_IN5_4 ( port0, port1, sel, portY );
  input [4:0] port0;
  input [4:0] port1;
  output [4:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, n1, n2, n3, n4, n5, n6, n8, n9;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;

  BUF_X1 U1 ( .A(sel), .Z(n1) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n2) );
  INV_X1 U3 ( .A(n5), .ZN(N3) );
  AOI22_X1 U4 ( .A1(port0[2]), .A2(n3), .B1(port1[2]), .B2(n1), .ZN(n6) );
  AOI22_X1 U5 ( .A1(port0[1]), .A2(n3), .B1(port1[1]), .B2(n1), .ZN(n5) );
  INV_X1 U6 ( .A(n6), .ZN(N4) );
  INV_X1 U7 ( .A(n4), .ZN(N2) );
  AOI22_X1 U8 ( .A1(port0[0]), .A2(n3), .B1(port1[0]), .B2(n1), .ZN(n4) );
  AOI22_X1 U9 ( .A1(port0[4]), .A2(n3), .B1(n2), .B2(port1[4]), .ZN(n9) );
  INV_X1 U10 ( .A(n9), .ZN(N6) );
  AOI22_X1 U11 ( .A1(port0[3]), .A2(n3), .B1(port1[3]), .B2(n1), .ZN(n8) );
  INV_X1 U12 ( .A(n8), .ZN(N5) );
  INV_X1 U13 ( .A(n2), .ZN(n3) );
endmodule


module Mux_NBit_2x1_NBIT_IN5_2 ( port0, port1, sel, portY );
  input [4:0] port0;
  input [4:0] port1;
  output [4:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, n1, n2, n3, n4, n5, n6;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;

  INV_X1 U1 ( .A(sel), .ZN(n5) );
  INV_X1 U2 ( .A(n3), .ZN(N4) );
  AOI22_X1 U3 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(sel), .ZN(n3) );
  INV_X1 U4 ( .A(n2), .ZN(N3) );
  AOI22_X1 U5 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(sel), .ZN(n2) );
  INV_X1 U6 ( .A(n4), .ZN(N5) );
  AOI22_X1 U7 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(sel), .ZN(n4) );
  INV_X1 U8 ( .A(n1), .ZN(N2) );
  AOI22_X1 U9 ( .A1(port0[0]), .A2(n5), .B1(port1[0]), .B2(sel), .ZN(n1) );
  INV_X1 U10 ( .A(n6), .ZN(N6) );
  AOI22_X1 U11 ( .A1(port0[4]), .A2(n5), .B1(sel), .B2(port1[4]), .ZN(n6) );
endmodule


module Mux_NBit_2x1_NBIT_IN5_1 ( port0, port1, sel, portY );
  input [4:0] port0;
  input [4:0] port1;
  output [4:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, n1, n2, n3, n4, n5, n6;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;

  INV_X1 U1 ( .A(sel), .ZN(n5) );
  INV_X1 U2 ( .A(n1), .ZN(N2) );
  AOI22_X1 U3 ( .A1(port0[0]), .A2(n5), .B1(port1[0]), .B2(sel), .ZN(n1) );
  INV_X1 U4 ( .A(n2), .ZN(N3) );
  AOI22_X1 U5 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(sel), .ZN(n2) );
  INV_X1 U6 ( .A(n3), .ZN(N4) );
  AOI22_X1 U7 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(sel), .ZN(n3) );
  INV_X1 U8 ( .A(n4), .ZN(N5) );
  AOI22_X1 U9 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(sel), .ZN(n4) );
  INV_X1 U10 ( .A(n6), .ZN(N6) );
  AOI22_X1 U11 ( .A1(port0[4]), .A2(n5), .B1(sel), .B2(port1[4]), .ZN(n6) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_120 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  INV_X1 U16 ( .A(n59), .ZN(N4) );
  INV_X1 U17 ( .A(n60), .ZN(N5) );
  INV_X1 U18 ( .A(n61), .ZN(N6) );
  INV_X1 U19 ( .A(n62), .ZN(N7) );
  INV_X1 U20 ( .A(n63), .ZN(N8) );
  INV_X1 U21 ( .A(n57), .ZN(N32) );
  INV_X1 U22 ( .A(n58), .ZN(N33) );
  INV_X1 U23 ( .A(n28), .ZN(N2) );
  INV_X1 U24 ( .A(n54), .ZN(N3) );
  INV_X1 U25 ( .A(n21), .ZN(N13) );
  INV_X1 U26 ( .A(n22), .ZN(N14) );
  INV_X1 U27 ( .A(n23), .ZN(N15) );
  INV_X1 U28 ( .A(n24), .ZN(N16) );
  INV_X1 U29 ( .A(n25), .ZN(N17) );
  INV_X1 U30 ( .A(n26), .ZN(N18) );
  INV_X1 U31 ( .A(n27), .ZN(N19) );
  INV_X1 U32 ( .A(n29), .ZN(N20) );
  INV_X1 U33 ( .A(n30), .ZN(N21) );
  INV_X1 U34 ( .A(n31), .ZN(N22) );
  INV_X1 U35 ( .A(n32), .ZN(N23) );
  INV_X1 U36 ( .A(n33), .ZN(N24) );
  INV_X1 U37 ( .A(n35), .ZN(N25) );
  INV_X1 U38 ( .A(n50), .ZN(N26) );
  INV_X1 U39 ( .A(n51), .ZN(N27) );
  INV_X1 U40 ( .A(n52), .ZN(N28) );
  INV_X1 U41 ( .A(n53), .ZN(N29) );
  INV_X1 U42 ( .A(n55), .ZN(N30) );
  INV_X1 U43 ( .A(n56), .ZN(N31) );
  INV_X1 U44 ( .A(n18), .ZN(N10) );
  INV_X1 U45 ( .A(n19), .ZN(N11) );
  INV_X1 U46 ( .A(n20), .ZN(N12) );
  AOI22_X1 U47 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U48 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U49 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U50 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U51 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U52 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U53 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U54 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U55 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U56 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U57 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U58 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U59 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U60 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U61 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U62 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U63 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U64 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U65 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U66 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_119 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  INV_X1 U16 ( .A(n59), .ZN(N4) );
  INV_X1 U17 ( .A(n60), .ZN(N5) );
  INV_X1 U18 ( .A(n61), .ZN(N6) );
  INV_X1 U19 ( .A(n62), .ZN(N7) );
  INV_X1 U20 ( .A(n63), .ZN(N8) );
  INV_X1 U21 ( .A(n57), .ZN(N32) );
  INV_X1 U22 ( .A(n58), .ZN(N33) );
  INV_X1 U23 ( .A(n28), .ZN(N2) );
  INV_X1 U24 ( .A(n54), .ZN(N3) );
  INV_X1 U25 ( .A(n21), .ZN(N13) );
  INV_X1 U26 ( .A(n22), .ZN(N14) );
  INV_X1 U27 ( .A(n23), .ZN(N15) );
  INV_X1 U28 ( .A(n24), .ZN(N16) );
  INV_X1 U29 ( .A(n25), .ZN(N17) );
  INV_X1 U30 ( .A(n26), .ZN(N18) );
  INV_X1 U31 ( .A(n27), .ZN(N19) );
  INV_X1 U32 ( .A(n29), .ZN(N20) );
  INV_X1 U33 ( .A(n30), .ZN(N21) );
  INV_X1 U34 ( .A(n31), .ZN(N22) );
  INV_X1 U35 ( .A(n32), .ZN(N23) );
  INV_X1 U36 ( .A(n33), .ZN(N24) );
  INV_X1 U37 ( .A(n35), .ZN(N25) );
  INV_X1 U38 ( .A(n50), .ZN(N26) );
  INV_X1 U39 ( .A(n51), .ZN(N27) );
  INV_X1 U40 ( .A(n52), .ZN(N28) );
  INV_X1 U41 ( .A(n53), .ZN(N29) );
  INV_X1 U42 ( .A(n55), .ZN(N30) );
  INV_X1 U43 ( .A(n56), .ZN(N31) );
  INV_X1 U44 ( .A(n18), .ZN(N10) );
  INV_X1 U45 ( .A(n19), .ZN(N11) );
  INV_X1 U46 ( .A(n20), .ZN(N12) );
  AOI22_X1 U47 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U48 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U49 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U50 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U51 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U52 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U53 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U54 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U55 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U56 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U57 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U58 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U59 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U60 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U61 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U62 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U63 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U64 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U65 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U66 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_118 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  INV_X1 U16 ( .A(n59), .ZN(N4) );
  INV_X1 U17 ( .A(n60), .ZN(N5) );
  INV_X1 U18 ( .A(n61), .ZN(N6) );
  INV_X1 U19 ( .A(n62), .ZN(N7) );
  INV_X1 U20 ( .A(n63), .ZN(N8) );
  INV_X1 U21 ( .A(n57), .ZN(N32) );
  INV_X1 U22 ( .A(n58), .ZN(N33) );
  INV_X1 U23 ( .A(n28), .ZN(N2) );
  INV_X1 U24 ( .A(n54), .ZN(N3) );
  INV_X1 U25 ( .A(n21), .ZN(N13) );
  INV_X1 U26 ( .A(n22), .ZN(N14) );
  INV_X1 U27 ( .A(n23), .ZN(N15) );
  INV_X1 U28 ( .A(n24), .ZN(N16) );
  INV_X1 U29 ( .A(n25), .ZN(N17) );
  INV_X1 U30 ( .A(n26), .ZN(N18) );
  INV_X1 U31 ( .A(n27), .ZN(N19) );
  INV_X1 U32 ( .A(n29), .ZN(N20) );
  INV_X1 U33 ( .A(n30), .ZN(N21) );
  INV_X1 U34 ( .A(n31), .ZN(N22) );
  INV_X1 U35 ( .A(n32), .ZN(N23) );
  INV_X1 U36 ( .A(n33), .ZN(N24) );
  INV_X1 U37 ( .A(n35), .ZN(N25) );
  INV_X1 U38 ( .A(n50), .ZN(N26) );
  INV_X1 U39 ( .A(n51), .ZN(N27) );
  INV_X1 U40 ( .A(n52), .ZN(N28) );
  INV_X1 U41 ( .A(n53), .ZN(N29) );
  INV_X1 U42 ( .A(n55), .ZN(N30) );
  INV_X1 U43 ( .A(n56), .ZN(N31) );
  INV_X1 U44 ( .A(n18), .ZN(N10) );
  INV_X1 U45 ( .A(n19), .ZN(N11) );
  INV_X1 U46 ( .A(n20), .ZN(N12) );
  AOI22_X1 U47 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U48 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U49 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U50 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U51 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U52 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U53 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U54 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U55 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U56 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U57 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U58 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U59 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U60 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U61 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U62 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U63 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U64 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U65 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U66 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_117 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n59), .ZN(N4) );
  AOI22_X1 U16 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U17 ( .A(n60), .ZN(N5) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U19 ( .A(n61), .ZN(N6) );
  AOI22_X1 U20 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U21 ( .A(n62), .ZN(N7) );
  AOI22_X1 U22 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U23 ( .A(n63), .ZN(N8) );
  AOI22_X1 U24 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U25 ( .A(n64), .ZN(N9) );
  AOI22_X1 U26 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U31 ( .A(n28), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U33 ( .A(n54), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U35 ( .A(n18), .ZN(N10) );
  AOI22_X1 U36 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U37 ( .A(n19), .ZN(N11) );
  AOI22_X1 U38 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U39 ( .A(n20), .ZN(N12) );
  AOI22_X1 U40 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U41 ( .A(n21), .ZN(N13) );
  AOI22_X1 U42 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U43 ( .A(n22), .ZN(N14) );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U45 ( .A(n23), .ZN(N15) );
  AOI22_X1 U46 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U47 ( .A(n24), .ZN(N16) );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U49 ( .A(n25), .ZN(N17) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U51 ( .A(n26), .ZN(N18) );
  AOI22_X1 U52 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U53 ( .A(n27), .ZN(N19) );
  AOI22_X1 U54 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U55 ( .A(n29), .ZN(N20) );
  AOI22_X1 U56 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U57 ( .A(n30), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U59 ( .A(n31), .ZN(N22) );
  AOI22_X1 U60 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U61 ( .A(n32), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U63 ( .A(n33), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U65 ( .A(n35), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U67 ( .A(n50), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U69 ( .A(n51), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U71 ( .A(n52), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U73 ( .A(n53), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U75 ( .A(n55), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_116 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  AOI22_X1 U18 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U19 ( .A(n60), .ZN(N5) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U21 ( .A(n61), .ZN(N6) );
  AOI22_X1 U22 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U23 ( .A(n62), .ZN(N7) );
  AOI22_X1 U24 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U25 ( .A(n63), .ZN(N8) );
  AOI22_X1 U26 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U31 ( .A(n28), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U33 ( .A(n54), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U35 ( .A(n18), .ZN(N10) );
  AOI22_X1 U36 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U37 ( .A(n19), .ZN(N11) );
  AOI22_X1 U38 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U39 ( .A(n20), .ZN(N12) );
  AOI22_X1 U40 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U41 ( .A(n21), .ZN(N13) );
  AOI22_X1 U42 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U43 ( .A(n22), .ZN(N14) );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U45 ( .A(n23), .ZN(N15) );
  AOI22_X1 U46 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U47 ( .A(n24), .ZN(N16) );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U49 ( .A(n25), .ZN(N17) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U51 ( .A(n26), .ZN(N18) );
  AOI22_X1 U52 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U53 ( .A(n27), .ZN(N19) );
  AOI22_X1 U54 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U55 ( .A(n29), .ZN(N20) );
  AOI22_X1 U56 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U57 ( .A(n30), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U59 ( .A(n31), .ZN(N22) );
  AOI22_X1 U60 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U61 ( .A(n32), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U63 ( .A(n33), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U65 ( .A(n35), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U67 ( .A(n50), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U69 ( .A(n51), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U71 ( .A(n52), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U73 ( .A(n53), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U75 ( .A(n55), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_115 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n59), .ZN(N4) );
  AOI22_X1 U16 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U17 ( .A(n60), .ZN(N5) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U19 ( .A(n61), .ZN(N6) );
  AOI22_X1 U20 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U21 ( .A(n62), .ZN(N7) );
  AOI22_X1 U22 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U23 ( .A(n63), .ZN(N8) );
  AOI22_X1 U24 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U25 ( .A(n57), .ZN(N32) );
  AOI22_X1 U26 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U27 ( .A(n58), .ZN(N33) );
  AOI22_X1 U28 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U29 ( .A(n28), .ZN(N2) );
  AOI22_X1 U30 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U31 ( .A(n54), .ZN(N3) );
  AOI22_X1 U32 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U33 ( .A(n18), .ZN(N10) );
  AOI22_X1 U34 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U35 ( .A(n19), .ZN(N11) );
  AOI22_X1 U36 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U37 ( .A(n20), .ZN(N12) );
  AOI22_X1 U38 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U39 ( .A(n21), .ZN(N13) );
  AOI22_X1 U40 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U41 ( .A(n22), .ZN(N14) );
  AOI22_X1 U42 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U43 ( .A(n23), .ZN(N15) );
  AOI22_X1 U44 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U45 ( .A(n24), .ZN(N16) );
  AOI22_X1 U46 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U47 ( .A(n25), .ZN(N17) );
  AOI22_X1 U48 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U49 ( .A(n26), .ZN(N18) );
  AOI22_X1 U50 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U51 ( .A(n27), .ZN(N19) );
  AOI22_X1 U52 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U53 ( .A(n29), .ZN(N20) );
  AOI22_X1 U54 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U55 ( .A(n30), .ZN(N21) );
  AOI22_X1 U56 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U57 ( .A(n31), .ZN(N22) );
  AOI22_X1 U58 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U59 ( .A(n32), .ZN(N23) );
  AOI22_X1 U60 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U61 ( .A(n33), .ZN(N24) );
  AOI22_X1 U62 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U63 ( .A(n35), .ZN(N25) );
  AOI22_X1 U64 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U65 ( .A(n50), .ZN(N26) );
  AOI22_X1 U66 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U67 ( .A(n51), .ZN(N27) );
  AOI22_X1 U68 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U69 ( .A(n52), .ZN(N28) );
  AOI22_X1 U70 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U71 ( .A(n53), .ZN(N29) );
  AOI22_X1 U72 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U73 ( .A(n55), .ZN(N30) );
  AOI22_X1 U74 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U75 ( .A(n56), .ZN(N31) );
  AOI22_X1 U76 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U77 ( .A(n64), .ZN(N9) );
  AOI22_X1 U78 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_114 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  AOI22_X1 U15 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U16 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U17 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U18 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U19 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U20 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U21 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U22 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U23 ( .A(n59), .ZN(N4) );
  INV_X1 U24 ( .A(n60), .ZN(N5) );
  INV_X1 U25 ( .A(n61), .ZN(N6) );
  INV_X1 U26 ( .A(n62), .ZN(N7) );
  INV_X1 U27 ( .A(n63), .ZN(N8) );
  INV_X1 U28 ( .A(n57), .ZN(N32) );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U31 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U32 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U33 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U34 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U35 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U36 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U37 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U38 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U39 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U40 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U41 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U42 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U43 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U44 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U45 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U46 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U47 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U48 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U49 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U50 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U51 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U52 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U53 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U54 ( .A(n28), .ZN(N2) );
  INV_X1 U55 ( .A(n54), .ZN(N3) );
  INV_X1 U56 ( .A(n18), .ZN(N10) );
  INV_X1 U57 ( .A(n19), .ZN(N11) );
  INV_X1 U58 ( .A(n20), .ZN(N12) );
  INV_X1 U59 ( .A(n21), .ZN(N13) );
  INV_X1 U60 ( .A(n22), .ZN(N14) );
  INV_X1 U61 ( .A(n23), .ZN(N15) );
  INV_X1 U62 ( .A(n24), .ZN(N16) );
  INV_X1 U63 ( .A(n25), .ZN(N17) );
  INV_X1 U64 ( .A(n26), .ZN(N18) );
  INV_X1 U65 ( .A(n27), .ZN(N19) );
  INV_X1 U66 ( .A(n29), .ZN(N20) );
  INV_X1 U67 ( .A(n30), .ZN(N21) );
  INV_X1 U68 ( .A(n31), .ZN(N22) );
  INV_X1 U69 ( .A(n32), .ZN(N23) );
  INV_X1 U70 ( .A(n33), .ZN(N24) );
  INV_X1 U71 ( .A(n35), .ZN(N25) );
  INV_X1 U72 ( .A(n50), .ZN(N26) );
  INV_X1 U73 ( .A(n51), .ZN(N27) );
  INV_X1 U74 ( .A(n52), .ZN(N28) );
  INV_X1 U75 ( .A(n53), .ZN(N29) );
  INV_X1 U76 ( .A(n55), .ZN(N30) );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  INV_X1 U78 ( .A(n64), .ZN(N9) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_113 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  AOI22_X1 U18 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U19 ( .A(n60), .ZN(N5) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U21 ( .A(n61), .ZN(N6) );
  AOI22_X1 U22 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U23 ( .A(n62), .ZN(N7) );
  AOI22_X1 U24 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U25 ( .A(n63), .ZN(N8) );
  AOI22_X1 U26 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U31 ( .A(n28), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U33 ( .A(n54), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U35 ( .A(n18), .ZN(N10) );
  AOI22_X1 U36 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U37 ( .A(n19), .ZN(N11) );
  AOI22_X1 U38 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U39 ( .A(n20), .ZN(N12) );
  AOI22_X1 U40 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U41 ( .A(n21), .ZN(N13) );
  AOI22_X1 U42 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U43 ( .A(n22), .ZN(N14) );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U45 ( .A(n23), .ZN(N15) );
  AOI22_X1 U46 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U47 ( .A(n24), .ZN(N16) );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U49 ( .A(n25), .ZN(N17) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U51 ( .A(n26), .ZN(N18) );
  AOI22_X1 U52 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U53 ( .A(n27), .ZN(N19) );
  AOI22_X1 U54 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U55 ( .A(n29), .ZN(N20) );
  AOI22_X1 U56 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U57 ( .A(n30), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U59 ( .A(n31), .ZN(N22) );
  AOI22_X1 U60 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U61 ( .A(n32), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U63 ( .A(n33), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U65 ( .A(n35), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U67 ( .A(n50), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U69 ( .A(n51), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U71 ( .A(n52), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U73 ( .A(n53), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U75 ( .A(n55), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_112 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  AOI22_X1 U18 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U19 ( .A(n60), .ZN(N5) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U21 ( .A(n61), .ZN(N6) );
  AOI22_X1 U22 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U23 ( .A(n62), .ZN(N7) );
  AOI22_X1 U24 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U25 ( .A(n63), .ZN(N8) );
  AOI22_X1 U26 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U31 ( .A(n28), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U33 ( .A(n54), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U35 ( .A(n18), .ZN(N10) );
  AOI22_X1 U36 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U37 ( .A(n19), .ZN(N11) );
  AOI22_X1 U38 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U39 ( .A(n20), .ZN(N12) );
  AOI22_X1 U40 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U41 ( .A(n21), .ZN(N13) );
  AOI22_X1 U42 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U43 ( .A(n22), .ZN(N14) );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U45 ( .A(n23), .ZN(N15) );
  AOI22_X1 U46 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U47 ( .A(n24), .ZN(N16) );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U49 ( .A(n25), .ZN(N17) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U51 ( .A(n26), .ZN(N18) );
  AOI22_X1 U52 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U53 ( .A(n27), .ZN(N19) );
  AOI22_X1 U54 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U55 ( .A(n29), .ZN(N20) );
  AOI22_X1 U56 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U57 ( .A(n30), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U59 ( .A(n31), .ZN(N22) );
  AOI22_X1 U60 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U61 ( .A(n32), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U63 ( .A(n33), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U65 ( .A(n35), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U67 ( .A(n50), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U69 ( .A(n51), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U71 ( .A(n52), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U73 ( .A(n53), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U75 ( .A(n55), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_111 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  AOI22_X1 U18 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U19 ( .A(n60), .ZN(N5) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U21 ( .A(n61), .ZN(N6) );
  AOI22_X1 U22 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U23 ( .A(n62), .ZN(N7) );
  AOI22_X1 U24 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U25 ( .A(n63), .ZN(N8) );
  AOI22_X1 U26 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U31 ( .A(n28), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U33 ( .A(n54), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U35 ( .A(n18), .ZN(N10) );
  AOI22_X1 U36 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U37 ( .A(n19), .ZN(N11) );
  AOI22_X1 U38 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U39 ( .A(n20), .ZN(N12) );
  AOI22_X1 U40 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U41 ( .A(n21), .ZN(N13) );
  AOI22_X1 U42 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U43 ( .A(n22), .ZN(N14) );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U45 ( .A(n23), .ZN(N15) );
  AOI22_X1 U46 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U47 ( .A(n24), .ZN(N16) );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U49 ( .A(n25), .ZN(N17) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U51 ( .A(n26), .ZN(N18) );
  AOI22_X1 U52 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U53 ( .A(n27), .ZN(N19) );
  AOI22_X1 U54 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U55 ( .A(n29), .ZN(N20) );
  AOI22_X1 U56 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U57 ( .A(n30), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U59 ( .A(n31), .ZN(N22) );
  AOI22_X1 U60 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U61 ( .A(n32), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U63 ( .A(n33), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U65 ( .A(n35), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U67 ( .A(n50), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U69 ( .A(n51), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U71 ( .A(n52), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U73 ( .A(n53), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U75 ( .A(n55), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_110 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U17 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U18 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U19 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U20 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U21 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U22 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U23 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U24 ( .A(n59), .ZN(N4) );
  INV_X1 U25 ( .A(n60), .ZN(N5) );
  INV_X1 U26 ( .A(n61), .ZN(N6) );
  INV_X1 U27 ( .A(n62), .ZN(N7) );
  INV_X1 U28 ( .A(n63), .ZN(N8) );
  INV_X1 U29 ( .A(n57), .ZN(N32) );
  INV_X1 U30 ( .A(n58), .ZN(N33) );
  AOI22_X1 U31 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U32 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U33 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U34 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U35 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U36 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U37 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U38 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U39 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U40 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U41 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U42 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U43 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U44 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U45 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U46 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U47 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U48 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U49 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U50 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U51 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U52 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U53 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U54 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U55 ( .A(n28), .ZN(N2) );
  INV_X1 U56 ( .A(n54), .ZN(N3) );
  INV_X1 U57 ( .A(n18), .ZN(N10) );
  INV_X1 U58 ( .A(n19), .ZN(N11) );
  INV_X1 U59 ( .A(n20), .ZN(N12) );
  INV_X1 U60 ( .A(n21), .ZN(N13) );
  INV_X1 U61 ( .A(n22), .ZN(N14) );
  INV_X1 U62 ( .A(n23), .ZN(N15) );
  INV_X1 U63 ( .A(n24), .ZN(N16) );
  INV_X1 U64 ( .A(n25), .ZN(N17) );
  INV_X1 U65 ( .A(n26), .ZN(N18) );
  INV_X1 U66 ( .A(n27), .ZN(N19) );
  INV_X1 U67 ( .A(n29), .ZN(N20) );
  INV_X1 U68 ( .A(n30), .ZN(N21) );
  INV_X1 U69 ( .A(n31), .ZN(N22) );
  INV_X1 U70 ( .A(n32), .ZN(N23) );
  INV_X1 U71 ( .A(n33), .ZN(N24) );
  INV_X1 U72 ( .A(n35), .ZN(N25) );
  INV_X1 U73 ( .A(n50), .ZN(N26) );
  INV_X1 U74 ( .A(n51), .ZN(N27) );
  INV_X1 U75 ( .A(n52), .ZN(N28) );
  INV_X1 U76 ( .A(n53), .ZN(N29) );
  INV_X1 U77 ( .A(n55), .ZN(N30) );
  INV_X1 U78 ( .A(n56), .ZN(N31) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_109 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n59), .ZN(N4) );
  INV_X1 U16 ( .A(n60), .ZN(N5) );
  INV_X1 U17 ( .A(n61), .ZN(N6) );
  INV_X1 U18 ( .A(n62), .ZN(N7) );
  INV_X1 U19 ( .A(n63), .ZN(N8) );
  INV_X1 U20 ( .A(n57), .ZN(N32) );
  INV_X1 U21 ( .A(n58), .ZN(N33) );
  INV_X1 U22 ( .A(n28), .ZN(N2) );
  INV_X1 U23 ( .A(n54), .ZN(N3) );
  INV_X1 U24 ( .A(n21), .ZN(N13) );
  INV_X1 U25 ( .A(n22), .ZN(N14) );
  INV_X1 U26 ( .A(n23), .ZN(N15) );
  INV_X1 U27 ( .A(n24), .ZN(N16) );
  INV_X1 U28 ( .A(n25), .ZN(N17) );
  INV_X1 U29 ( .A(n26), .ZN(N18) );
  INV_X1 U30 ( .A(n27), .ZN(N19) );
  INV_X1 U31 ( .A(n29), .ZN(N20) );
  INV_X1 U32 ( .A(n30), .ZN(N21) );
  INV_X1 U33 ( .A(n31), .ZN(N22) );
  INV_X1 U34 ( .A(n32), .ZN(N23) );
  INV_X1 U35 ( .A(n33), .ZN(N24) );
  INV_X1 U36 ( .A(n35), .ZN(N25) );
  INV_X1 U37 ( .A(n50), .ZN(N26) );
  INV_X1 U38 ( .A(n51), .ZN(N27) );
  INV_X1 U39 ( .A(n52), .ZN(N28) );
  INV_X1 U40 ( .A(n53), .ZN(N29) );
  INV_X1 U41 ( .A(n55), .ZN(N30) );
  INV_X1 U42 ( .A(n56), .ZN(N31) );
  INV_X1 U43 ( .A(n18), .ZN(N10) );
  INV_X1 U44 ( .A(n19), .ZN(N11) );
  INV_X1 U45 ( .A(n20), .ZN(N12) );
  AOI22_X1 U46 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U47 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U48 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U49 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U50 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U51 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U52 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U53 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U54 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U55 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U56 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U57 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U58 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U59 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U60 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U61 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U62 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U63 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U64 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U65 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U66 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U67 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U68 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U69 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U70 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U71 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U72 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U73 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U75 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U76 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U77 ( .A(n64), .ZN(N9) );
  AOI22_X1 U78 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_108 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n59), .ZN(N4) );
  INV_X1 U16 ( .A(n60), .ZN(N5) );
  INV_X1 U17 ( .A(n61), .ZN(N6) );
  INV_X1 U18 ( .A(n62), .ZN(N7) );
  INV_X1 U19 ( .A(n63), .ZN(N8) );
  INV_X1 U20 ( .A(n57), .ZN(N32) );
  INV_X1 U21 ( .A(n58), .ZN(N33) );
  INV_X1 U22 ( .A(n28), .ZN(N2) );
  INV_X1 U23 ( .A(n54), .ZN(N3) );
  INV_X1 U24 ( .A(n21), .ZN(N13) );
  INV_X1 U25 ( .A(n22), .ZN(N14) );
  INV_X1 U26 ( .A(n23), .ZN(N15) );
  INV_X1 U27 ( .A(n24), .ZN(N16) );
  INV_X1 U28 ( .A(n25), .ZN(N17) );
  INV_X1 U29 ( .A(n26), .ZN(N18) );
  INV_X1 U30 ( .A(n27), .ZN(N19) );
  INV_X1 U31 ( .A(n29), .ZN(N20) );
  INV_X1 U32 ( .A(n30), .ZN(N21) );
  INV_X1 U33 ( .A(n31), .ZN(N22) );
  INV_X1 U34 ( .A(n32), .ZN(N23) );
  INV_X1 U35 ( .A(n33), .ZN(N24) );
  INV_X1 U36 ( .A(n35), .ZN(N25) );
  INV_X1 U37 ( .A(n50), .ZN(N26) );
  INV_X1 U38 ( .A(n51), .ZN(N27) );
  INV_X1 U39 ( .A(n52), .ZN(N28) );
  INV_X1 U40 ( .A(n53), .ZN(N29) );
  INV_X1 U41 ( .A(n55), .ZN(N30) );
  INV_X1 U42 ( .A(n56), .ZN(N31) );
  INV_X1 U43 ( .A(n18), .ZN(N10) );
  INV_X1 U44 ( .A(n19), .ZN(N11) );
  INV_X1 U45 ( .A(n20), .ZN(N12) );
  AOI22_X1 U46 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U47 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U48 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U49 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U50 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U51 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U52 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U53 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U54 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U55 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U56 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U57 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U58 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U59 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U60 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U61 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U62 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U63 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U64 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U65 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U66 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U67 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U68 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U69 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U70 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U71 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U72 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U73 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U75 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U76 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U77 ( .A(n64), .ZN(N9) );
  AOI22_X1 U78 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_107 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n59), .ZN(N4) );
  INV_X1 U16 ( .A(n60), .ZN(N5) );
  INV_X1 U17 ( .A(n61), .ZN(N6) );
  INV_X1 U18 ( .A(n62), .ZN(N7) );
  INV_X1 U19 ( .A(n63), .ZN(N8) );
  INV_X1 U20 ( .A(n57), .ZN(N32) );
  INV_X1 U21 ( .A(n58), .ZN(N33) );
  INV_X1 U22 ( .A(n28), .ZN(N2) );
  INV_X1 U23 ( .A(n54), .ZN(N3) );
  INV_X1 U24 ( .A(n21), .ZN(N13) );
  INV_X1 U25 ( .A(n22), .ZN(N14) );
  INV_X1 U26 ( .A(n23), .ZN(N15) );
  INV_X1 U27 ( .A(n24), .ZN(N16) );
  INV_X1 U28 ( .A(n25), .ZN(N17) );
  INV_X1 U29 ( .A(n26), .ZN(N18) );
  INV_X1 U30 ( .A(n27), .ZN(N19) );
  INV_X1 U31 ( .A(n29), .ZN(N20) );
  INV_X1 U32 ( .A(n30), .ZN(N21) );
  INV_X1 U33 ( .A(n31), .ZN(N22) );
  INV_X1 U34 ( .A(n32), .ZN(N23) );
  INV_X1 U35 ( .A(n33), .ZN(N24) );
  INV_X1 U36 ( .A(n35), .ZN(N25) );
  INV_X1 U37 ( .A(n50), .ZN(N26) );
  INV_X1 U38 ( .A(n51), .ZN(N27) );
  INV_X1 U39 ( .A(n52), .ZN(N28) );
  INV_X1 U40 ( .A(n53), .ZN(N29) );
  INV_X1 U41 ( .A(n55), .ZN(N30) );
  INV_X1 U42 ( .A(n56), .ZN(N31) );
  INV_X1 U43 ( .A(n18), .ZN(N10) );
  INV_X1 U44 ( .A(n19), .ZN(N11) );
  INV_X1 U45 ( .A(n20), .ZN(N12) );
  AOI22_X1 U46 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U47 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U48 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U49 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U50 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U51 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U52 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U53 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U54 ( .A(n64), .ZN(N9) );
  AOI22_X1 U55 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U56 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U57 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U58 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U59 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U60 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U61 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U62 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U63 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U64 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U65 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U66 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_106 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  INV_X1 U12 ( .A(n59), .ZN(N4) );
  INV_X1 U13 ( .A(n60), .ZN(N5) );
  INV_X1 U14 ( .A(n61), .ZN(N6) );
  INV_X1 U15 ( .A(n62), .ZN(N7) );
  INV_X1 U16 ( .A(n63), .ZN(N8) );
  INV_X1 U17 ( .A(n57), .ZN(N32) );
  INV_X1 U18 ( .A(n58), .ZN(N33) );
  BUF_X1 U19 ( .A(sel), .Z(n6) );
  BUF_X1 U20 ( .A(sel), .Z(n5) );
  BUF_X1 U21 ( .A(sel), .Z(n4) );
  INV_X1 U22 ( .A(n28), .ZN(N2) );
  INV_X1 U23 ( .A(n54), .ZN(N3) );
  INV_X1 U24 ( .A(n21), .ZN(N13) );
  INV_X1 U25 ( .A(n22), .ZN(N14) );
  INV_X1 U26 ( .A(n23), .ZN(N15) );
  INV_X1 U27 ( .A(n24), .ZN(N16) );
  INV_X1 U28 ( .A(n25), .ZN(N17) );
  INV_X1 U29 ( .A(n26), .ZN(N18) );
  INV_X1 U30 ( .A(n27), .ZN(N19) );
  INV_X1 U31 ( .A(n29), .ZN(N20) );
  INV_X1 U32 ( .A(n30), .ZN(N21) );
  INV_X1 U33 ( .A(n31), .ZN(N22) );
  INV_X1 U34 ( .A(n32), .ZN(N23) );
  INV_X1 U35 ( .A(n33), .ZN(N24) );
  INV_X1 U36 ( .A(n35), .ZN(N25) );
  INV_X1 U37 ( .A(n50), .ZN(N26) );
  INV_X1 U38 ( .A(n51), .ZN(N27) );
  INV_X1 U39 ( .A(n52), .ZN(N28) );
  INV_X1 U40 ( .A(n53), .ZN(N29) );
  INV_X1 U41 ( .A(n55), .ZN(N30) );
  INV_X1 U42 ( .A(n56), .ZN(N31) );
  INV_X1 U43 ( .A(n18), .ZN(N10) );
  INV_X1 U44 ( .A(n19), .ZN(N11) );
  INV_X1 U45 ( .A(n20), .ZN(N12) );
  AOI22_X1 U46 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U47 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U48 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U49 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U50 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U51 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U52 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U53 ( .A(n64), .ZN(N9) );
  AOI22_X1 U54 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U55 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U56 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U57 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U58 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U59 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U60 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U61 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U62 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U63 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U64 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U65 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U66 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_105 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  INV_X1 U12 ( .A(n64), .ZN(N9) );
  AOI22_X1 U13 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U14 ( .A(n59), .ZN(N4) );
  AOI22_X1 U15 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U16 ( .A(n60), .ZN(N5) );
  AOI22_X1 U17 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U18 ( .A(n61), .ZN(N6) );
  AOI22_X1 U19 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U20 ( .A(n62), .ZN(N7) );
  AOI22_X1 U21 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U22 ( .A(n63), .ZN(N8) );
  AOI22_X1 U23 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U24 ( .A(n57), .ZN(N32) );
  AOI22_X1 U25 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U26 ( .A(n58), .ZN(N33) );
  AOI22_X1 U27 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U28 ( .A(n28), .ZN(N2) );
  AOI22_X1 U29 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U30 ( .A(n54), .ZN(N3) );
  AOI22_X1 U31 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U32 ( .A(n21), .ZN(N13) );
  AOI22_X1 U33 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U34 ( .A(n22), .ZN(N14) );
  AOI22_X1 U35 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U36 ( .A(n23), .ZN(N15) );
  AOI22_X1 U37 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U38 ( .A(n24), .ZN(N16) );
  AOI22_X1 U39 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U40 ( .A(n25), .ZN(N17) );
  AOI22_X1 U41 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U42 ( .A(n26), .ZN(N18) );
  AOI22_X1 U43 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U44 ( .A(n27), .ZN(N19) );
  AOI22_X1 U45 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U46 ( .A(n29), .ZN(N20) );
  AOI22_X1 U47 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U48 ( .A(n30), .ZN(N21) );
  AOI22_X1 U49 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U50 ( .A(n31), .ZN(N22) );
  AOI22_X1 U51 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U52 ( .A(n32), .ZN(N23) );
  AOI22_X1 U53 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U54 ( .A(n33), .ZN(N24) );
  AOI22_X1 U55 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U56 ( .A(n35), .ZN(N25) );
  AOI22_X1 U57 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U58 ( .A(n50), .ZN(N26) );
  AOI22_X1 U59 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U60 ( .A(n51), .ZN(N27) );
  AOI22_X1 U61 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U62 ( .A(n52), .ZN(N28) );
  AOI22_X1 U63 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U64 ( .A(n53), .ZN(N29) );
  AOI22_X1 U65 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U66 ( .A(n55), .ZN(N30) );
  AOI22_X1 U67 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U68 ( .A(n56), .ZN(N31) );
  AOI22_X1 U69 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U70 ( .A(n18), .ZN(N10) );
  AOI22_X1 U71 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U72 ( .A(n19), .ZN(N11) );
  AOI22_X1 U73 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U74 ( .A(n20), .ZN(N12) );
  AOI22_X1 U75 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  BUF_X1 U76 ( .A(sel), .Z(n6) );
  BUF_X1 U77 ( .A(sel), .Z(n5) );
  BUF_X1 U78 ( .A(sel), .Z(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_104 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  INV_X1 U12 ( .A(n64), .ZN(N9) );
  AOI22_X1 U13 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U14 ( .A(n59), .ZN(N4) );
  AOI22_X1 U15 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U16 ( .A(n60), .ZN(N5) );
  AOI22_X1 U17 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U18 ( .A(n61), .ZN(N6) );
  AOI22_X1 U19 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U20 ( .A(n62), .ZN(N7) );
  AOI22_X1 U21 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U22 ( .A(n63), .ZN(N8) );
  AOI22_X1 U23 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U24 ( .A(n57), .ZN(N32) );
  AOI22_X1 U25 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U26 ( .A(n58), .ZN(N33) );
  AOI22_X1 U27 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U28 ( .A(n28), .ZN(N2) );
  AOI22_X1 U29 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U30 ( .A(n54), .ZN(N3) );
  AOI22_X1 U31 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U32 ( .A(n21), .ZN(N13) );
  AOI22_X1 U33 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U34 ( .A(n22), .ZN(N14) );
  AOI22_X1 U35 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U36 ( .A(n23), .ZN(N15) );
  AOI22_X1 U37 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U38 ( .A(n24), .ZN(N16) );
  AOI22_X1 U39 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U40 ( .A(n25), .ZN(N17) );
  AOI22_X1 U41 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U42 ( .A(n26), .ZN(N18) );
  AOI22_X1 U43 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U44 ( .A(n27), .ZN(N19) );
  AOI22_X1 U45 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U46 ( .A(n29), .ZN(N20) );
  AOI22_X1 U47 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U48 ( .A(n30), .ZN(N21) );
  AOI22_X1 U49 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U50 ( .A(n31), .ZN(N22) );
  AOI22_X1 U51 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U52 ( .A(n32), .ZN(N23) );
  AOI22_X1 U53 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U54 ( .A(n33), .ZN(N24) );
  AOI22_X1 U55 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U56 ( .A(n35), .ZN(N25) );
  AOI22_X1 U57 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U58 ( .A(n50), .ZN(N26) );
  AOI22_X1 U59 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U60 ( .A(n51), .ZN(N27) );
  AOI22_X1 U61 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U62 ( .A(n52), .ZN(N28) );
  AOI22_X1 U63 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U64 ( .A(n53), .ZN(N29) );
  AOI22_X1 U65 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U66 ( .A(n55), .ZN(N30) );
  AOI22_X1 U67 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U68 ( .A(n56), .ZN(N31) );
  AOI22_X1 U69 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U70 ( .A(n18), .ZN(N10) );
  AOI22_X1 U71 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U72 ( .A(n19), .ZN(N11) );
  AOI22_X1 U73 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U74 ( .A(n20), .ZN(N12) );
  AOI22_X1 U75 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  BUF_X1 U76 ( .A(sel), .Z(n6) );
  BUF_X1 U77 ( .A(sel), .Z(n5) );
  BUF_X1 U78 ( .A(sel), .Z(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_103 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  INV_X1 U12 ( .A(n59), .ZN(N4) );
  AOI22_X1 U13 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U14 ( .A(n60), .ZN(N5) );
  AOI22_X1 U15 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U16 ( .A(n61), .ZN(N6) );
  AOI22_X1 U17 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U18 ( .A(n62), .ZN(N7) );
  AOI22_X1 U19 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U20 ( .A(n63), .ZN(N8) );
  AOI22_X1 U21 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U22 ( .A(n57), .ZN(N32) );
  AOI22_X1 U23 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U24 ( .A(n58), .ZN(N33) );
  AOI22_X1 U25 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U26 ( .A(n28), .ZN(N2) );
  AOI22_X1 U27 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U28 ( .A(n54), .ZN(N3) );
  AOI22_X1 U29 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U30 ( .A(n18), .ZN(N10) );
  AOI22_X1 U31 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U32 ( .A(n19), .ZN(N11) );
  AOI22_X1 U33 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U34 ( .A(n20), .ZN(N12) );
  AOI22_X1 U35 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U36 ( .A(n21), .ZN(N13) );
  AOI22_X1 U37 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U38 ( .A(n22), .ZN(N14) );
  AOI22_X1 U39 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U40 ( .A(n23), .ZN(N15) );
  AOI22_X1 U41 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U42 ( .A(n24), .ZN(N16) );
  AOI22_X1 U43 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U44 ( .A(n25), .ZN(N17) );
  AOI22_X1 U45 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U46 ( .A(n26), .ZN(N18) );
  AOI22_X1 U47 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U48 ( .A(n27), .ZN(N19) );
  AOI22_X1 U49 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U50 ( .A(n29), .ZN(N20) );
  AOI22_X1 U51 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U52 ( .A(n30), .ZN(N21) );
  AOI22_X1 U53 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U54 ( .A(n31), .ZN(N22) );
  AOI22_X1 U55 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U56 ( .A(n32), .ZN(N23) );
  AOI22_X1 U57 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U58 ( .A(n33), .ZN(N24) );
  AOI22_X1 U59 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U60 ( .A(n35), .ZN(N25) );
  AOI22_X1 U61 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U62 ( .A(n50), .ZN(N26) );
  AOI22_X1 U63 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U64 ( .A(n51), .ZN(N27) );
  AOI22_X1 U65 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U66 ( .A(n52), .ZN(N28) );
  AOI22_X1 U67 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U68 ( .A(n53), .ZN(N29) );
  AOI22_X1 U69 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U70 ( .A(n55), .ZN(N30) );
  AOI22_X1 U71 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U72 ( .A(n56), .ZN(N31) );
  AOI22_X1 U73 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U74 ( .A(n64), .ZN(N9) );
  AOI22_X1 U75 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  BUF_X1 U76 ( .A(sel), .Z(n6) );
  BUF_X1 U77 ( .A(sel), .Z(n5) );
  BUF_X1 U78 ( .A(sel), .Z(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_102 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  INV_X1 U12 ( .A(n59), .ZN(N4) );
  INV_X1 U13 ( .A(n60), .ZN(N5) );
  INV_X1 U14 ( .A(n61), .ZN(N6) );
  INV_X1 U15 ( .A(n62), .ZN(N7) );
  INV_X1 U16 ( .A(n63), .ZN(N8) );
  INV_X1 U17 ( .A(n57), .ZN(N32) );
  INV_X1 U18 ( .A(n58), .ZN(N33) );
  INV_X1 U19 ( .A(n28), .ZN(N2) );
  INV_X1 U20 ( .A(n54), .ZN(N3) );
  INV_X1 U21 ( .A(n18), .ZN(N10) );
  INV_X1 U22 ( .A(n19), .ZN(N11) );
  INV_X1 U23 ( .A(n20), .ZN(N12) );
  INV_X1 U24 ( .A(n21), .ZN(N13) );
  INV_X1 U25 ( .A(n22), .ZN(N14) );
  INV_X1 U26 ( .A(n23), .ZN(N15) );
  INV_X1 U27 ( .A(n24), .ZN(N16) );
  INV_X1 U28 ( .A(n25), .ZN(N17) );
  INV_X1 U29 ( .A(n26), .ZN(N18) );
  INV_X1 U30 ( .A(n27), .ZN(N19) );
  INV_X1 U31 ( .A(n29), .ZN(N20) );
  INV_X1 U32 ( .A(n30), .ZN(N21) );
  INV_X1 U33 ( .A(n31), .ZN(N22) );
  INV_X1 U34 ( .A(n32), .ZN(N23) );
  INV_X1 U35 ( .A(n33), .ZN(N24) );
  INV_X1 U36 ( .A(n35), .ZN(N25) );
  INV_X1 U37 ( .A(n50), .ZN(N26) );
  INV_X1 U38 ( .A(n51), .ZN(N27) );
  INV_X1 U39 ( .A(n52), .ZN(N28) );
  INV_X1 U40 ( .A(n53), .ZN(N29) );
  INV_X1 U41 ( .A(n55), .ZN(N30) );
  INV_X1 U42 ( .A(n56), .ZN(N31) );
  INV_X1 U43 ( .A(n64), .ZN(N9) );
  BUF_X1 U44 ( .A(sel), .Z(n6) );
  BUF_X1 U45 ( .A(sel), .Z(n5) );
  BUF_X1 U46 ( .A(sel), .Z(n4) );
  AOI22_X1 U47 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U48 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U49 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U50 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U51 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U52 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U53 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U54 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U55 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U56 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U57 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U58 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U59 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U60 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U61 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U62 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U63 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U64 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U65 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U66 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U67 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U68 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U69 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U70 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U71 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U72 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U73 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U74 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U75 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U77 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  AOI22_X1 U78 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_101 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  INV_X1 U12 ( .A(n59), .ZN(N4) );
  AOI22_X1 U13 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U14 ( .A(n60), .ZN(N5) );
  AOI22_X1 U15 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U16 ( .A(n61), .ZN(N6) );
  AOI22_X1 U17 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U18 ( .A(n62), .ZN(N7) );
  AOI22_X1 U19 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U20 ( .A(n63), .ZN(N8) );
  AOI22_X1 U21 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U22 ( .A(n57), .ZN(N32) );
  AOI22_X1 U23 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U24 ( .A(n58), .ZN(N33) );
  AOI22_X1 U25 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U26 ( .A(n28), .ZN(N2) );
  AOI22_X1 U27 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U28 ( .A(n54), .ZN(N3) );
  AOI22_X1 U29 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U30 ( .A(n18), .ZN(N10) );
  AOI22_X1 U31 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U32 ( .A(n19), .ZN(N11) );
  AOI22_X1 U33 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U34 ( .A(n20), .ZN(N12) );
  AOI22_X1 U35 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U36 ( .A(n21), .ZN(N13) );
  AOI22_X1 U37 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U38 ( .A(n22), .ZN(N14) );
  AOI22_X1 U39 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U40 ( .A(n23), .ZN(N15) );
  AOI22_X1 U41 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U42 ( .A(n24), .ZN(N16) );
  AOI22_X1 U43 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U44 ( .A(n25), .ZN(N17) );
  AOI22_X1 U45 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U46 ( .A(n26), .ZN(N18) );
  AOI22_X1 U47 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U48 ( .A(n27), .ZN(N19) );
  AOI22_X1 U49 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U50 ( .A(n29), .ZN(N20) );
  AOI22_X1 U51 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U52 ( .A(n30), .ZN(N21) );
  AOI22_X1 U53 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U54 ( .A(n31), .ZN(N22) );
  AOI22_X1 U55 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U56 ( .A(n32), .ZN(N23) );
  AOI22_X1 U57 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U58 ( .A(n33), .ZN(N24) );
  AOI22_X1 U59 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U60 ( .A(n35), .ZN(N25) );
  AOI22_X1 U61 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U62 ( .A(n50), .ZN(N26) );
  AOI22_X1 U63 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U64 ( .A(n51), .ZN(N27) );
  AOI22_X1 U65 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U66 ( .A(n52), .ZN(N28) );
  AOI22_X1 U67 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U68 ( .A(n53), .ZN(N29) );
  AOI22_X1 U69 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U70 ( .A(n55), .ZN(N30) );
  AOI22_X1 U71 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U72 ( .A(n56), .ZN(N31) );
  AOI22_X1 U73 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U74 ( .A(n64), .ZN(N9) );
  AOI22_X1 U75 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  BUF_X1 U76 ( .A(sel), .Z(n6) );
  BUF_X1 U77 ( .A(sel), .Z(n5) );
  BUF_X1 U78 ( .A(sel), .Z(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_100 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  INV_X1 U12 ( .A(n59), .ZN(N4) );
  INV_X1 U13 ( .A(n60), .ZN(N5) );
  INV_X1 U14 ( .A(n61), .ZN(N6) );
  INV_X1 U15 ( .A(n62), .ZN(N7) );
  INV_X1 U16 ( .A(n63), .ZN(N8) );
  INV_X1 U17 ( .A(n57), .ZN(N32) );
  INV_X1 U18 ( .A(n58), .ZN(N33) );
  INV_X1 U19 ( .A(n28), .ZN(N2) );
  INV_X1 U20 ( .A(n54), .ZN(N3) );
  INV_X1 U21 ( .A(n18), .ZN(N10) );
  INV_X1 U22 ( .A(n19), .ZN(N11) );
  INV_X1 U23 ( .A(n20), .ZN(N12) );
  INV_X1 U24 ( .A(n21), .ZN(N13) );
  INV_X1 U25 ( .A(n22), .ZN(N14) );
  INV_X1 U26 ( .A(n23), .ZN(N15) );
  INV_X1 U27 ( .A(n24), .ZN(N16) );
  INV_X1 U28 ( .A(n25), .ZN(N17) );
  INV_X1 U29 ( .A(n26), .ZN(N18) );
  INV_X1 U30 ( .A(n27), .ZN(N19) );
  INV_X1 U31 ( .A(n29), .ZN(N20) );
  INV_X1 U32 ( .A(n30), .ZN(N21) );
  INV_X1 U33 ( .A(n31), .ZN(N22) );
  INV_X1 U34 ( .A(n32), .ZN(N23) );
  INV_X1 U35 ( .A(n33), .ZN(N24) );
  INV_X1 U36 ( .A(n35), .ZN(N25) );
  INV_X1 U37 ( .A(n50), .ZN(N26) );
  INV_X1 U38 ( .A(n51), .ZN(N27) );
  INV_X1 U39 ( .A(n52), .ZN(N28) );
  INV_X1 U40 ( .A(n53), .ZN(N29) );
  INV_X1 U41 ( .A(n55), .ZN(N30) );
  INV_X1 U42 ( .A(n56), .ZN(N31) );
  INV_X1 U43 ( .A(n64), .ZN(N9) );
  AOI22_X1 U44 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  BUF_X1 U45 ( .A(sel), .Z(n6) );
  BUF_X1 U46 ( .A(sel), .Z(n5) );
  BUF_X1 U47 ( .A(sel), .Z(n4) );
  AOI22_X1 U48 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U49 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U50 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U51 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U52 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U53 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U54 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U55 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U56 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U57 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U58 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U59 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U60 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U61 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U62 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U63 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U64 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U65 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U66 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_99 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  INV_X1 U12 ( .A(n64), .ZN(N9) );
  AOI22_X1 U13 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U14 ( .A(n59), .ZN(N4) );
  AOI22_X1 U15 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U16 ( .A(n60), .ZN(N5) );
  AOI22_X1 U17 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U18 ( .A(n61), .ZN(N6) );
  AOI22_X1 U19 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U20 ( .A(n62), .ZN(N7) );
  AOI22_X1 U21 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U22 ( .A(n63), .ZN(N8) );
  AOI22_X1 U23 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U24 ( .A(n57), .ZN(N32) );
  AOI22_X1 U25 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U26 ( .A(n58), .ZN(N33) );
  AOI22_X1 U27 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U28 ( .A(n28), .ZN(N2) );
  AOI22_X1 U29 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U30 ( .A(n54), .ZN(N3) );
  AOI22_X1 U31 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U32 ( .A(n21), .ZN(N13) );
  AOI22_X1 U33 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U34 ( .A(n22), .ZN(N14) );
  AOI22_X1 U35 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U36 ( .A(n23), .ZN(N15) );
  AOI22_X1 U37 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U38 ( .A(n24), .ZN(N16) );
  AOI22_X1 U39 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U40 ( .A(n25), .ZN(N17) );
  AOI22_X1 U41 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U42 ( .A(n26), .ZN(N18) );
  AOI22_X1 U43 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U44 ( .A(n27), .ZN(N19) );
  AOI22_X1 U45 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U46 ( .A(n29), .ZN(N20) );
  AOI22_X1 U47 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U48 ( .A(n30), .ZN(N21) );
  AOI22_X1 U49 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U50 ( .A(n31), .ZN(N22) );
  AOI22_X1 U51 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U52 ( .A(n32), .ZN(N23) );
  AOI22_X1 U53 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U54 ( .A(n33), .ZN(N24) );
  AOI22_X1 U55 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U56 ( .A(n35), .ZN(N25) );
  AOI22_X1 U57 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U58 ( .A(n50), .ZN(N26) );
  AOI22_X1 U59 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U60 ( .A(n51), .ZN(N27) );
  AOI22_X1 U61 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U62 ( .A(n52), .ZN(N28) );
  AOI22_X1 U63 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U64 ( .A(n53), .ZN(N29) );
  AOI22_X1 U65 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U66 ( .A(n55), .ZN(N30) );
  AOI22_X1 U67 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U68 ( .A(n56), .ZN(N31) );
  AOI22_X1 U69 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U70 ( .A(n18), .ZN(N10) );
  AOI22_X1 U71 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U72 ( .A(n19), .ZN(N11) );
  AOI22_X1 U73 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U74 ( .A(n20), .ZN(N12) );
  AOI22_X1 U75 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  BUF_X1 U76 ( .A(sel), .Z(n6) );
  BUF_X1 U77 ( .A(sel), .Z(n5) );
  BUF_X1 U78 ( .A(sel), .Z(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_98 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  INV_X1 U12 ( .A(n64), .ZN(N9) );
  INV_X1 U13 ( .A(n59), .ZN(N4) );
  AOI22_X1 U14 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U15 ( .A(n60), .ZN(N5) );
  AOI22_X1 U16 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U17 ( .A(n61), .ZN(N6) );
  AOI22_X1 U18 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U19 ( .A(n62), .ZN(N7) );
  AOI22_X1 U20 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U21 ( .A(n63), .ZN(N8) );
  AOI22_X1 U22 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U23 ( .A(n57), .ZN(N32) );
  AOI22_X1 U24 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U25 ( .A(n58), .ZN(N33) );
  AOI22_X1 U26 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U27 ( .A(n28), .ZN(N2) );
  AOI22_X1 U28 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U29 ( .A(n54), .ZN(N3) );
  AOI22_X1 U30 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U31 ( .A(n21), .ZN(N13) );
  AOI22_X1 U32 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U33 ( .A(n22), .ZN(N14) );
  AOI22_X1 U34 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U35 ( .A(n23), .ZN(N15) );
  AOI22_X1 U36 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U37 ( .A(n24), .ZN(N16) );
  AOI22_X1 U38 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U39 ( .A(n25), .ZN(N17) );
  AOI22_X1 U40 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U41 ( .A(n26), .ZN(N18) );
  AOI22_X1 U42 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U43 ( .A(n27), .ZN(N19) );
  AOI22_X1 U44 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U45 ( .A(n29), .ZN(N20) );
  AOI22_X1 U46 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U47 ( .A(n30), .ZN(N21) );
  AOI22_X1 U48 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U49 ( .A(n31), .ZN(N22) );
  AOI22_X1 U50 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U51 ( .A(n32), .ZN(N23) );
  AOI22_X1 U52 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U53 ( .A(n33), .ZN(N24) );
  AOI22_X1 U54 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U55 ( .A(n35), .ZN(N25) );
  AOI22_X1 U56 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U57 ( .A(n50), .ZN(N26) );
  AOI22_X1 U58 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U59 ( .A(n51), .ZN(N27) );
  AOI22_X1 U60 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U61 ( .A(n52), .ZN(N28) );
  AOI22_X1 U62 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U63 ( .A(n53), .ZN(N29) );
  AOI22_X1 U64 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U65 ( .A(n55), .ZN(N30) );
  AOI22_X1 U66 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U67 ( .A(n56), .ZN(N31) );
  AOI22_X1 U68 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U69 ( .A(n18), .ZN(N10) );
  AOI22_X1 U70 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U71 ( .A(n19), .ZN(N11) );
  AOI22_X1 U72 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U73 ( .A(n20), .ZN(N12) );
  AOI22_X1 U74 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  BUF_X1 U75 ( .A(sel), .Z(n6) );
  BUF_X1 U76 ( .A(sel), .Z(n5) );
  BUF_X1 U77 ( .A(sel), .Z(n4) );
  AOI22_X1 U78 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_97 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  INV_X1 U3 ( .A(n59), .ZN(N4) );
  AOI22_X1 U4 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U5 ( .A(n60), .ZN(N5) );
  AOI22_X1 U6 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U7 ( .A(n61), .ZN(N6) );
  AOI22_X1 U8 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U9 ( .A(n62), .ZN(N7) );
  AOI22_X1 U10 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U11 ( .A(n63), .ZN(N8) );
  AOI22_X1 U12 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U13 ( .A(n57), .ZN(N32) );
  AOI22_X1 U14 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U15 ( .A(n58), .ZN(N33) );
  AOI22_X1 U16 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U17 ( .A(n28), .ZN(N2) );
  AOI22_X1 U18 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U19 ( .A(n54), .ZN(N3) );
  AOI22_X1 U20 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U21 ( .A(n18), .ZN(N10) );
  AOI22_X1 U22 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U23 ( .A(n19), .ZN(N11) );
  AOI22_X1 U24 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U25 ( .A(n20), .ZN(N12) );
  AOI22_X1 U26 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U27 ( .A(n21), .ZN(N13) );
  AOI22_X1 U28 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U29 ( .A(n22), .ZN(N14) );
  AOI22_X1 U30 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U31 ( .A(n23), .ZN(N15) );
  AOI22_X1 U32 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U33 ( .A(n24), .ZN(N16) );
  AOI22_X1 U34 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U35 ( .A(n25), .ZN(N17) );
  AOI22_X1 U36 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U37 ( .A(n26), .ZN(N18) );
  AOI22_X1 U38 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U39 ( .A(n27), .ZN(N19) );
  AOI22_X1 U40 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U41 ( .A(n29), .ZN(N20) );
  AOI22_X1 U42 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U43 ( .A(n30), .ZN(N21) );
  AOI22_X1 U44 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U45 ( .A(n31), .ZN(N22) );
  AOI22_X1 U46 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U47 ( .A(n32), .ZN(N23) );
  AOI22_X1 U48 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U49 ( .A(n33), .ZN(N24) );
  AOI22_X1 U50 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U51 ( .A(n35), .ZN(N25) );
  AOI22_X1 U52 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U53 ( .A(n50), .ZN(N26) );
  AOI22_X1 U54 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U55 ( .A(n51), .ZN(N27) );
  AOI22_X1 U56 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U57 ( .A(n52), .ZN(N28) );
  AOI22_X1 U58 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U59 ( .A(n53), .ZN(N29) );
  AOI22_X1 U60 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U61 ( .A(n55), .ZN(N30) );
  AOI22_X1 U62 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U63 ( .A(n56), .ZN(N31) );
  AOI22_X1 U64 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U65 ( .A(n64), .ZN(N9) );
  AOI22_X1 U66 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  BUF_X1 U67 ( .A(n4), .Z(n9) );
  BUF_X1 U68 ( .A(n6), .Z(n15) );
  BUF_X1 U69 ( .A(n5), .Z(n14) );
  BUF_X1 U70 ( .A(n5), .Z(n12) );
  BUF_X1 U71 ( .A(n4), .Z(n11) );
  BUF_X1 U72 ( .A(n5), .Z(n13) );
  BUF_X1 U73 ( .A(n4), .Z(n10) );
  BUF_X1 U74 ( .A(n6), .Z(n17) );
  BUF_X1 U75 ( .A(n6), .Z(n16) );
  BUF_X1 U76 ( .A(sel), .Z(n6) );
  BUF_X1 U77 ( .A(sel), .Z(n5) );
  BUF_X1 U78 ( .A(sel), .Z(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_96 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  INV_X1 U3 ( .A(n59), .ZN(N4) );
  INV_X1 U4 ( .A(n60), .ZN(N5) );
  INV_X1 U5 ( .A(n61), .ZN(N6) );
  INV_X1 U6 ( .A(n62), .ZN(N7) );
  INV_X1 U7 ( .A(n63), .ZN(N8) );
  INV_X1 U8 ( .A(n57), .ZN(N32) );
  INV_X1 U9 ( .A(n58), .ZN(N33) );
  INV_X1 U10 ( .A(n28), .ZN(N2) );
  INV_X1 U11 ( .A(n54), .ZN(N3) );
  INV_X1 U12 ( .A(n18), .ZN(N10) );
  INV_X1 U13 ( .A(n19), .ZN(N11) );
  INV_X1 U14 ( .A(n20), .ZN(N12) );
  INV_X1 U15 ( .A(n21), .ZN(N13) );
  INV_X1 U16 ( .A(n22), .ZN(N14) );
  INV_X1 U17 ( .A(n23), .ZN(N15) );
  INV_X1 U18 ( .A(n24), .ZN(N16) );
  INV_X1 U19 ( .A(n25), .ZN(N17) );
  INV_X1 U20 ( .A(n26), .ZN(N18) );
  INV_X1 U21 ( .A(n27), .ZN(N19) );
  INV_X1 U22 ( .A(n29), .ZN(N20) );
  INV_X1 U23 ( .A(n30), .ZN(N21) );
  INV_X1 U24 ( .A(n31), .ZN(N22) );
  INV_X1 U25 ( .A(n32), .ZN(N23) );
  INV_X1 U26 ( .A(n33), .ZN(N24) );
  INV_X1 U27 ( .A(n35), .ZN(N25) );
  INV_X1 U28 ( .A(n50), .ZN(N26) );
  INV_X1 U29 ( .A(n51), .ZN(N27) );
  INV_X1 U30 ( .A(n52), .ZN(N28) );
  INV_X1 U31 ( .A(n53), .ZN(N29) );
  INV_X1 U32 ( .A(n55), .ZN(N30) );
  INV_X1 U33 ( .A(n56), .ZN(N31) );
  INV_X1 U34 ( .A(n64), .ZN(N9) );
  BUF_X1 U35 ( .A(n4), .Z(n9) );
  BUF_X1 U36 ( .A(n6), .Z(n15) );
  BUF_X1 U37 ( .A(n5), .Z(n14) );
  BUF_X1 U38 ( .A(n5), .Z(n12) );
  BUF_X1 U39 ( .A(n4), .Z(n11) );
  BUF_X1 U40 ( .A(n5), .Z(n13) );
  BUF_X1 U41 ( .A(n4), .Z(n10) );
  BUF_X1 U42 ( .A(n6), .Z(n17) );
  BUF_X1 U43 ( .A(n6), .Z(n16) );
  AOI22_X1 U44 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U45 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U46 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U47 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U48 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U49 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U50 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U51 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U52 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U53 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U54 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U55 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U56 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U57 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U58 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U59 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U60 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U61 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U62 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U63 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U64 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U65 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U66 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U67 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U68 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U69 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U71 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U72 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U73 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U74 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  AOI22_X1 U75 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  BUF_X1 U76 ( .A(sel), .Z(n6) );
  BUF_X1 U77 ( .A(sel), .Z(n5) );
  BUF_X1 U78 ( .A(sel), .Z(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_95 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  INV_X1 U3 ( .A(n59), .ZN(N4) );
  INV_X1 U4 ( .A(n60), .ZN(N5) );
  INV_X1 U5 ( .A(n61), .ZN(N6) );
  INV_X1 U6 ( .A(n62), .ZN(N7) );
  INV_X1 U7 ( .A(n63), .ZN(N8) );
  INV_X1 U8 ( .A(n57), .ZN(N32) );
  INV_X1 U9 ( .A(n58), .ZN(N33) );
  INV_X1 U10 ( .A(n28), .ZN(N2) );
  INV_X1 U11 ( .A(n54), .ZN(N3) );
  INV_X1 U12 ( .A(n18), .ZN(N10) );
  INV_X1 U13 ( .A(n19), .ZN(N11) );
  INV_X1 U14 ( .A(n20), .ZN(N12) );
  INV_X1 U15 ( .A(n21), .ZN(N13) );
  INV_X1 U16 ( .A(n22), .ZN(N14) );
  INV_X1 U17 ( .A(n23), .ZN(N15) );
  INV_X1 U18 ( .A(n24), .ZN(N16) );
  INV_X1 U19 ( .A(n25), .ZN(N17) );
  INV_X1 U20 ( .A(n26), .ZN(N18) );
  INV_X1 U21 ( .A(n27), .ZN(N19) );
  INV_X1 U22 ( .A(n29), .ZN(N20) );
  INV_X1 U23 ( .A(n30), .ZN(N21) );
  INV_X1 U24 ( .A(n31), .ZN(N22) );
  INV_X1 U25 ( .A(n32), .ZN(N23) );
  INV_X1 U26 ( .A(n33), .ZN(N24) );
  INV_X1 U27 ( .A(n35), .ZN(N25) );
  INV_X1 U28 ( .A(n50), .ZN(N26) );
  INV_X1 U29 ( .A(n51), .ZN(N27) );
  INV_X1 U30 ( .A(n52), .ZN(N28) );
  INV_X1 U31 ( .A(n53), .ZN(N29) );
  INV_X1 U32 ( .A(n55), .ZN(N30) );
  INV_X1 U33 ( .A(n56), .ZN(N31) );
  INV_X1 U34 ( .A(n64), .ZN(N9) );
  AOI22_X1 U35 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  BUF_X1 U36 ( .A(n4), .Z(n9) );
  BUF_X1 U37 ( .A(n6), .Z(n15) );
  BUF_X1 U38 ( .A(n5), .Z(n14) );
  BUF_X1 U39 ( .A(n5), .Z(n12) );
  BUF_X1 U40 ( .A(n4), .Z(n11) );
  BUF_X1 U41 ( .A(n5), .Z(n13) );
  BUF_X1 U42 ( .A(n4), .Z(n10) );
  BUF_X1 U43 ( .A(n6), .Z(n17) );
  BUF_X1 U44 ( .A(n6), .Z(n16) );
  AOI22_X1 U45 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U46 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U47 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U48 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U49 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U50 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U51 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U52 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U53 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U54 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U55 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U56 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U57 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U58 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U59 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U60 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U61 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U62 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U63 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U64 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U65 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U66 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U67 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U68 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U69 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U70 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U71 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U73 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U74 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U75 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  BUF_X1 U76 ( .A(sel), .Z(n6) );
  BUF_X1 U77 ( .A(sel), .Z(n5) );
  BUF_X1 U78 ( .A(sel), .Z(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_94 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  INV_X1 U3 ( .A(n59), .ZN(N4) );
  AOI22_X1 U4 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U5 ( .A(n60), .ZN(N5) );
  AOI22_X1 U6 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U7 ( .A(n61), .ZN(N6) );
  AOI22_X1 U8 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U9 ( .A(n62), .ZN(N7) );
  AOI22_X1 U10 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U11 ( .A(n63), .ZN(N8) );
  AOI22_X1 U12 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U13 ( .A(n57), .ZN(N32) );
  AOI22_X1 U14 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U15 ( .A(n58), .ZN(N33) );
  AOI22_X1 U16 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U17 ( .A(n28), .ZN(N2) );
  AOI22_X1 U18 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U19 ( .A(n54), .ZN(N3) );
  AOI22_X1 U20 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U21 ( .A(n18), .ZN(N10) );
  AOI22_X1 U22 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U23 ( .A(n19), .ZN(N11) );
  AOI22_X1 U24 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U25 ( .A(n20), .ZN(N12) );
  AOI22_X1 U26 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U27 ( .A(n21), .ZN(N13) );
  AOI22_X1 U28 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U29 ( .A(n22), .ZN(N14) );
  AOI22_X1 U30 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U31 ( .A(n23), .ZN(N15) );
  AOI22_X1 U32 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U33 ( .A(n24), .ZN(N16) );
  AOI22_X1 U34 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U35 ( .A(n25), .ZN(N17) );
  AOI22_X1 U36 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U37 ( .A(n26), .ZN(N18) );
  AOI22_X1 U38 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U39 ( .A(n27), .ZN(N19) );
  AOI22_X1 U40 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U41 ( .A(n29), .ZN(N20) );
  AOI22_X1 U42 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U43 ( .A(n30), .ZN(N21) );
  AOI22_X1 U44 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U45 ( .A(n31), .ZN(N22) );
  AOI22_X1 U46 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U47 ( .A(n32), .ZN(N23) );
  AOI22_X1 U48 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U49 ( .A(n33), .ZN(N24) );
  AOI22_X1 U50 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U51 ( .A(n35), .ZN(N25) );
  AOI22_X1 U52 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U53 ( .A(n50), .ZN(N26) );
  AOI22_X1 U54 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U55 ( .A(n51), .ZN(N27) );
  AOI22_X1 U56 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U57 ( .A(n52), .ZN(N28) );
  AOI22_X1 U58 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U59 ( .A(n53), .ZN(N29) );
  AOI22_X1 U60 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U61 ( .A(n55), .ZN(N30) );
  AOI22_X1 U62 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U63 ( .A(n56), .ZN(N31) );
  AOI22_X1 U64 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U65 ( .A(n64), .ZN(N9) );
  BUF_X1 U66 ( .A(n4), .Z(n9) );
  BUF_X1 U67 ( .A(n6), .Z(n15) );
  BUF_X1 U68 ( .A(n5), .Z(n14) );
  BUF_X1 U69 ( .A(n5), .Z(n12) );
  BUF_X1 U70 ( .A(n4), .Z(n11) );
  BUF_X1 U71 ( .A(n5), .Z(n13) );
  BUF_X1 U72 ( .A(n4), .Z(n10) );
  BUF_X1 U73 ( .A(n6), .Z(n17) );
  BUF_X1 U74 ( .A(n6), .Z(n16) );
  AOI22_X1 U75 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  BUF_X1 U76 ( .A(sel), .Z(n6) );
  BUF_X1 U77 ( .A(sel), .Z(n5) );
  BUF_X1 U78 ( .A(sel), .Z(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_76 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n5), .Z(n14) );
  BUF_X1 U5 ( .A(n4), .Z(n11) );
  BUF_X1 U6 ( .A(n4), .Z(n10) );
  BUF_X1 U7 ( .A(n6), .Z(n17) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n61), .ZN(N6) );
  INV_X1 U16 ( .A(n60), .ZN(N5) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  INV_X1 U18 ( .A(n28), .ZN(N2) );
  INV_X1 U19 ( .A(n54), .ZN(N3) );
  INV_X1 U20 ( .A(n62), .ZN(N7) );
  INV_X1 U21 ( .A(n64), .ZN(N9) );
  INV_X1 U22 ( .A(n63), .ZN(N8) );
  INV_X1 U23 ( .A(n58), .ZN(N33) );
  INV_X1 U24 ( .A(n57), .ZN(N32) );
  INV_X1 U25 ( .A(n30), .ZN(N21) );
  INV_X1 U26 ( .A(n25), .ZN(N17) );
  INV_X1 U27 ( .A(n26), .ZN(N18) );
  INV_X1 U28 ( .A(n31), .ZN(N22) );
  INV_X1 U29 ( .A(n32), .ZN(N23) );
  INV_X1 U30 ( .A(n33), .ZN(N24) );
  INV_X1 U31 ( .A(n35), .ZN(N25) );
  INV_X1 U32 ( .A(n50), .ZN(N26) );
  INV_X1 U33 ( .A(n51), .ZN(N27) );
  INV_X1 U34 ( .A(n52), .ZN(N28) );
  INV_X1 U35 ( .A(n53), .ZN(N29) );
  INV_X1 U36 ( .A(n55), .ZN(N30) );
  INV_X1 U37 ( .A(n56), .ZN(N31) );
  INV_X1 U38 ( .A(n27), .ZN(N19) );
  INV_X1 U39 ( .A(n23), .ZN(N15) );
  INV_X1 U40 ( .A(n22), .ZN(N14) );
  INV_X1 U41 ( .A(n24), .ZN(N16) );
  INV_X1 U42 ( .A(n21), .ZN(N13) );
  INV_X1 U43 ( .A(n29), .ZN(N20) );
  INV_X1 U44 ( .A(n20), .ZN(N12) );
  INV_X1 U45 ( .A(n19), .ZN(N11) );
  INV_X1 U46 ( .A(n18), .ZN(N10) );
  AOI22_X1 U47 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U48 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U49 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U50 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U51 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U52 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U53 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U54 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U55 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U56 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U57 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U58 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U59 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U60 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U61 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U62 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U63 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U64 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U65 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U66 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_72 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n5), .Z(n14) );
  BUF_X1 U5 ( .A(n4), .Z(n11) );
  BUF_X1 U6 ( .A(n4), .Z(n10) );
  BUF_X1 U7 ( .A(n6), .Z(n17) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n61), .ZN(N6) );
  INV_X1 U16 ( .A(n60), .ZN(N5) );
  AOI22_X1 U17 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U18 ( .A(n59), .ZN(N4) );
  AOI22_X1 U19 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U21 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U22 ( .A(n28), .ZN(N2) );
  AOI22_X1 U23 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U24 ( .A(n54), .ZN(N3) );
  INV_X1 U25 ( .A(n62), .ZN(N7) );
  AOI22_X1 U26 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U27 ( .A(n64), .ZN(N9) );
  AOI22_X1 U28 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U29 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U30 ( .A(n63), .ZN(N8) );
  AOI22_X1 U31 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U32 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U33 ( .A(n58), .ZN(N33) );
  INV_X1 U34 ( .A(n57), .ZN(N32) );
  AOI22_X1 U35 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U36 ( .A(n29), .ZN(N20) );
  INV_X1 U37 ( .A(n27), .ZN(N19) );
  INV_X1 U38 ( .A(n20), .ZN(N12) );
  INV_X1 U39 ( .A(n23), .ZN(N15) );
  INV_X1 U40 ( .A(n22), .ZN(N14) );
  INV_X1 U41 ( .A(n24), .ZN(N16) );
  INV_X1 U42 ( .A(n19), .ZN(N11) );
  AOI22_X1 U43 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U44 ( .A(n18), .ZN(N10) );
  AOI22_X1 U45 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U46 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U47 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U48 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U49 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U51 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U52 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U53 ( .A(n21), .ZN(N13) );
  AOI22_X1 U54 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U55 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U56 ( .A(n30), .ZN(N21) );
  AOI22_X1 U57 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U58 ( .A(n31), .ZN(N22) );
  AOI22_X1 U59 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U60 ( .A(n32), .ZN(N23) );
  AOI22_X1 U61 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U62 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U63 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U64 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U65 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U66 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U67 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U68 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U69 ( .A(n25), .ZN(N17) );
  INV_X1 U70 ( .A(n26), .ZN(N18) );
  INV_X1 U71 ( .A(n33), .ZN(N24) );
  INV_X1 U72 ( .A(n35), .ZN(N25) );
  INV_X1 U73 ( .A(n50), .ZN(N26) );
  INV_X1 U74 ( .A(n51), .ZN(N27) );
  INV_X1 U75 ( .A(n52), .ZN(N28) );
  INV_X1 U76 ( .A(n53), .ZN(N29) );
  INV_X1 U77 ( .A(n55), .ZN(N30) );
  INV_X1 U78 ( .A(n56), .ZN(N31) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_68 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n5), .Z(n14) );
  BUF_X1 U5 ( .A(n4), .Z(n11) );
  BUF_X1 U6 ( .A(n4), .Z(n10) );
  BUF_X1 U7 ( .A(n6), .Z(n17) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n61), .ZN(N6) );
  INV_X1 U16 ( .A(n60), .ZN(N5) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  INV_X1 U18 ( .A(n54), .ZN(N3) );
  INV_X1 U19 ( .A(n62), .ZN(N7) );
  INV_X1 U20 ( .A(n58), .ZN(N33) );
  INV_X1 U21 ( .A(n57), .ZN(N32) );
  INV_X1 U22 ( .A(n24), .ZN(N16) );
  INV_X1 U23 ( .A(n21), .ZN(N13) );
  INV_X1 U24 ( .A(n30), .ZN(N21) );
  INV_X1 U25 ( .A(n31), .ZN(N22) );
  INV_X1 U26 ( .A(n32), .ZN(N23) );
  INV_X1 U27 ( .A(n64), .ZN(N9) );
  INV_X1 U28 ( .A(n63), .ZN(N8) );
  INV_X1 U29 ( .A(n25), .ZN(N17) );
  INV_X1 U30 ( .A(n26), .ZN(N18) );
  INV_X1 U31 ( .A(n33), .ZN(N24) );
  INV_X1 U32 ( .A(n35), .ZN(N25) );
  INV_X1 U33 ( .A(n50), .ZN(N26) );
  INV_X1 U34 ( .A(n51), .ZN(N27) );
  INV_X1 U35 ( .A(n52), .ZN(N28) );
  INV_X1 U36 ( .A(n53), .ZN(N29) );
  INV_X1 U37 ( .A(n55), .ZN(N30) );
  INV_X1 U38 ( .A(n56), .ZN(N31) );
  INV_X1 U39 ( .A(n29), .ZN(N20) );
  INV_X1 U40 ( .A(n27), .ZN(N19) );
  INV_X1 U41 ( .A(n23), .ZN(N15) );
  INV_X1 U42 ( .A(n22), .ZN(N14) );
  INV_X1 U43 ( .A(n20), .ZN(N12) );
  INV_X1 U44 ( .A(n19), .ZN(N11) );
  INV_X1 U45 ( .A(n18), .ZN(N10) );
  AOI22_X1 U46 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U47 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U48 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U49 ( .A(n28), .ZN(N2) );
  AOI22_X1 U50 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U51 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U52 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U53 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U54 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U55 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U56 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U57 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U58 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U59 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U60 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U61 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U62 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U63 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U64 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U65 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U66 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U67 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_63 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n5), .Z(n14) );
  BUF_X1 U4 ( .A(n4), .Z(n11) );
  BUF_X1 U5 ( .A(n4), .Z(n10) );
  BUF_X1 U6 ( .A(n6), .Z(n17) );
  BUF_X1 U7 ( .A(n4), .Z(n9) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n61), .ZN(N6) );
  AOI22_X1 U16 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U17 ( .A(n60), .ZN(N5) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U19 ( .A(n59), .ZN(N4) );
  AOI22_X1 U20 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U21 ( .A(n28), .ZN(N2) );
  AOI22_X1 U22 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U23 ( .A(n54), .ZN(N3) );
  AOI22_X1 U24 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U25 ( .A(n62), .ZN(N7) );
  AOI22_X1 U26 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U27 ( .A(n64), .ZN(N9) );
  AOI22_X1 U28 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U29 ( .A(n63), .ZN(N8) );
  AOI22_X1 U30 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U31 ( .A(n58), .ZN(N33) );
  AOI22_X1 U32 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U33 ( .A(n57), .ZN(N32) );
  AOI22_X1 U34 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U35 ( .A(n26), .ZN(N18) );
  AOI22_X1 U36 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U37 ( .A(n31), .ZN(N22) );
  AOI22_X1 U38 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U39 ( .A(n32), .ZN(N23) );
  AOI22_X1 U40 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U41 ( .A(n33), .ZN(N24) );
  AOI22_X1 U42 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U43 ( .A(n35), .ZN(N25) );
  AOI22_X1 U44 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U45 ( .A(n50), .ZN(N26) );
  AOI22_X1 U46 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U47 ( .A(n51), .ZN(N27) );
  AOI22_X1 U48 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U49 ( .A(n52), .ZN(N28) );
  AOI22_X1 U50 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U51 ( .A(n53), .ZN(N29) );
  AOI22_X1 U52 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U53 ( .A(n55), .ZN(N30) );
  AOI22_X1 U54 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U55 ( .A(n56), .ZN(N31) );
  AOI22_X1 U56 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U57 ( .A(n27), .ZN(N19) );
  AOI22_X1 U58 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U59 ( .A(n23), .ZN(N15) );
  AOI22_X1 U60 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U61 ( .A(n22), .ZN(N14) );
  AOI22_X1 U62 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U63 ( .A(n24), .ZN(N16) );
  AOI22_X1 U64 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U65 ( .A(n25), .ZN(N17) );
  AOI22_X1 U66 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U67 ( .A(n21), .ZN(N13) );
  AOI22_X1 U68 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U69 ( .A(n29), .ZN(N20) );
  AOI22_X1 U70 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U71 ( .A(n30), .ZN(N21) );
  AOI22_X1 U72 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U73 ( .A(n20), .ZN(N12) );
  AOI22_X1 U74 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U75 ( .A(n19), .ZN(N11) );
  AOI22_X1 U76 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U77 ( .A(n18), .ZN(N10) );
  AOI22_X1 U78 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_62 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n5), .Z(n14) );
  BUF_X1 U4 ( .A(n4), .Z(n11) );
  BUF_X1 U5 ( .A(n4), .Z(n10) );
  BUF_X1 U6 ( .A(n6), .Z(n17) );
  BUF_X1 U7 ( .A(n4), .Z(n9) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n61), .ZN(N6) );
  AOI22_X1 U16 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U17 ( .A(n60), .ZN(N5) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U19 ( .A(n59), .ZN(N4) );
  AOI22_X1 U20 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U21 ( .A(n28), .ZN(N2) );
  AOI22_X1 U22 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U23 ( .A(n54), .ZN(N3) );
  AOI22_X1 U24 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U25 ( .A(n62), .ZN(N7) );
  AOI22_X1 U26 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U27 ( .A(n64), .ZN(N9) );
  AOI22_X1 U28 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U29 ( .A(n63), .ZN(N8) );
  AOI22_X1 U30 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U31 ( .A(n58), .ZN(N33) );
  AOI22_X1 U32 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U33 ( .A(n57), .ZN(N32) );
  AOI22_X1 U34 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U35 ( .A(n30), .ZN(N21) );
  AOI22_X1 U36 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U37 ( .A(n25), .ZN(N17) );
  AOI22_X1 U38 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U39 ( .A(n26), .ZN(N18) );
  AOI22_X1 U40 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U41 ( .A(n31), .ZN(N22) );
  AOI22_X1 U42 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U43 ( .A(n32), .ZN(N23) );
  AOI22_X1 U44 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U45 ( .A(n33), .ZN(N24) );
  AOI22_X1 U46 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U47 ( .A(n35), .ZN(N25) );
  AOI22_X1 U48 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U49 ( .A(n50), .ZN(N26) );
  AOI22_X1 U50 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U51 ( .A(n51), .ZN(N27) );
  AOI22_X1 U52 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U53 ( .A(n52), .ZN(N28) );
  AOI22_X1 U54 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U55 ( .A(n53), .ZN(N29) );
  AOI22_X1 U56 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U57 ( .A(n55), .ZN(N30) );
  AOI22_X1 U58 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U59 ( .A(n56), .ZN(N31) );
  AOI22_X1 U60 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U61 ( .A(n27), .ZN(N19) );
  AOI22_X1 U62 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U63 ( .A(n23), .ZN(N15) );
  AOI22_X1 U64 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U65 ( .A(n22), .ZN(N14) );
  AOI22_X1 U66 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U67 ( .A(n24), .ZN(N16) );
  AOI22_X1 U68 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U69 ( .A(n21), .ZN(N13) );
  AOI22_X1 U70 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U71 ( .A(n29), .ZN(N20) );
  AOI22_X1 U72 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U73 ( .A(n20), .ZN(N12) );
  AOI22_X1 U74 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U75 ( .A(n19), .ZN(N11) );
  AOI22_X1 U76 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U77 ( .A(n18), .ZN(N10) );
  AOI22_X1 U78 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_61 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n8) );
  INV_X1 U2 ( .A(n17), .ZN(n7) );
  BUF_X1 U3 ( .A(n4), .Z(n11) );
  BUF_X1 U4 ( .A(n4), .Z(n10) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n6), .Z(n17) );
  BUF_X1 U7 ( .A(n4), .Z(n9) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n12) );
  BUF_X1 U11 ( .A(n5), .Z(n13) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n4) );
  BUF_X1 U14 ( .A(sel), .Z(n5) );
  INV_X1 U15 ( .A(n61), .ZN(N6) );
  AOI22_X1 U16 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U17 ( .A(n60), .ZN(N5) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U19 ( .A(n59), .ZN(N4) );
  AOI22_X1 U20 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U21 ( .A(n28), .ZN(N2) );
  AOI22_X1 U22 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U23 ( .A(n54), .ZN(N3) );
  AOI22_X1 U24 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U25 ( .A(n62), .ZN(N7) );
  AOI22_X1 U26 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U27 ( .A(n64), .ZN(N9) );
  AOI22_X1 U28 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U29 ( .A(n29), .ZN(N20) );
  AOI22_X1 U30 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U31 ( .A(n27), .ZN(N19) );
  AOI22_X1 U32 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U33 ( .A(n20), .ZN(N12) );
  AOI22_X1 U34 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U35 ( .A(n22), .ZN(N14) );
  AOI22_X1 U36 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U37 ( .A(n24), .ZN(N16) );
  AOI22_X1 U38 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U39 ( .A(n19), .ZN(N11) );
  AOI22_X1 U40 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U41 ( .A(n18), .ZN(N10) );
  AOI22_X1 U42 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U43 ( .A(n21), .ZN(N13) );
  AOI22_X1 U44 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U45 ( .A(n26), .ZN(N18) );
  AOI22_X1 U46 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U47 ( .A(n63), .ZN(N8) );
  AOI22_X1 U48 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U49 ( .A(n58), .ZN(N33) );
  AOI22_X1 U50 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U51 ( .A(n57), .ZN(N32) );
  AOI22_X1 U52 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U53 ( .A(n23), .ZN(N15) );
  AOI22_X1 U54 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U55 ( .A(n25), .ZN(N17) );
  AOI22_X1 U56 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U57 ( .A(n30), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U59 ( .A(n31), .ZN(N22) );
  AOI22_X1 U60 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U61 ( .A(n32), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U63 ( .A(n33), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U65 ( .A(n35), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U67 ( .A(n50), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U69 ( .A(n51), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U71 ( .A(n52), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U73 ( .A(n53), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U75 ( .A(n55), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_60 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n5), .Z(n14) );
  BUF_X1 U4 ( .A(n4), .Z(n11) );
  BUF_X1 U5 ( .A(n4), .Z(n10) );
  BUF_X1 U6 ( .A(n6), .Z(n17) );
  BUF_X1 U7 ( .A(n4), .Z(n9) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n61), .ZN(N6) );
  INV_X1 U16 ( .A(n60), .ZN(N5) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  INV_X1 U18 ( .A(n28), .ZN(N2) );
  INV_X1 U19 ( .A(n54), .ZN(N3) );
  INV_X1 U20 ( .A(n62), .ZN(N7) );
  INV_X1 U21 ( .A(n64), .ZN(N9) );
  INV_X1 U22 ( .A(n29), .ZN(N20) );
  INV_X1 U23 ( .A(n27), .ZN(N19) );
  INV_X1 U24 ( .A(n20), .ZN(N12) );
  INV_X1 U25 ( .A(n22), .ZN(N14) );
  INV_X1 U26 ( .A(n24), .ZN(N16) );
  INV_X1 U27 ( .A(n19), .ZN(N11) );
  INV_X1 U28 ( .A(n18), .ZN(N10) );
  INV_X1 U29 ( .A(n21), .ZN(N13) );
  INV_X1 U30 ( .A(n26), .ZN(N18) );
  INV_X1 U31 ( .A(n63), .ZN(N8) );
  INV_X1 U32 ( .A(n58), .ZN(N33) );
  INV_X1 U33 ( .A(n57), .ZN(N32) );
  INV_X1 U34 ( .A(n23), .ZN(N15) );
  INV_X1 U35 ( .A(n25), .ZN(N17) );
  INV_X1 U36 ( .A(n30), .ZN(N21) );
  INV_X1 U37 ( .A(n31), .ZN(N22) );
  INV_X1 U38 ( .A(n32), .ZN(N23) );
  INV_X1 U39 ( .A(n33), .ZN(N24) );
  INV_X1 U40 ( .A(n35), .ZN(N25) );
  INV_X1 U41 ( .A(n50), .ZN(N26) );
  INV_X1 U42 ( .A(n51), .ZN(N27) );
  INV_X1 U43 ( .A(n52), .ZN(N28) );
  INV_X1 U44 ( .A(n53), .ZN(N29) );
  INV_X1 U45 ( .A(n55), .ZN(N30) );
  INV_X1 U46 ( .A(n56), .ZN(N31) );
  AOI22_X1 U47 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U48 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U49 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U50 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U51 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U52 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U53 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U54 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U55 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U56 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U57 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U58 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U59 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U60 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U61 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U62 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U63 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U64 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U65 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U66 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U67 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U68 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U69 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U70 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_59 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n8) );
  INV_X1 U2 ( .A(n17), .ZN(n7) );
  BUF_X1 U3 ( .A(n4), .Z(n11) );
  BUF_X1 U4 ( .A(n4), .Z(n10) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n6), .Z(n17) );
  BUF_X1 U7 ( .A(n4), .Z(n9) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n28), .ZN(N2) );
  AOI22_X1 U16 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U17 ( .A(n61), .ZN(N6) );
  AOI22_X1 U18 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U19 ( .A(n60), .ZN(N5) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U21 ( .A(n59), .ZN(N4) );
  AOI22_X1 U22 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U23 ( .A(n54), .ZN(N3) );
  AOI22_X1 U24 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U25 ( .A(n62), .ZN(N7) );
  AOI22_X1 U26 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U27 ( .A(n64), .ZN(N9) );
  AOI22_X1 U28 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U29 ( .A(n63), .ZN(N8) );
  AOI22_X1 U30 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U31 ( .A(n58), .ZN(N33) );
  AOI22_X1 U32 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U33 ( .A(n57), .ZN(N32) );
  AOI22_X1 U34 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U35 ( .A(n22), .ZN(N14) );
  AOI22_X1 U36 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U37 ( .A(n26), .ZN(N18) );
  AOI22_X1 U38 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U39 ( .A(n31), .ZN(N22) );
  AOI22_X1 U40 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U41 ( .A(n32), .ZN(N23) );
  AOI22_X1 U42 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U43 ( .A(n33), .ZN(N24) );
  AOI22_X1 U44 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U45 ( .A(n35), .ZN(N25) );
  AOI22_X1 U46 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U47 ( .A(n50), .ZN(N26) );
  AOI22_X1 U48 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U49 ( .A(n51), .ZN(N27) );
  AOI22_X1 U50 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U51 ( .A(n52), .ZN(N28) );
  AOI22_X1 U52 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U53 ( .A(n53), .ZN(N29) );
  AOI22_X1 U54 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U55 ( .A(n55), .ZN(N30) );
  AOI22_X1 U56 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U57 ( .A(n56), .ZN(N31) );
  AOI22_X1 U58 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U59 ( .A(n27), .ZN(N19) );
  AOI22_X1 U60 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U61 ( .A(n23), .ZN(N15) );
  AOI22_X1 U62 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U63 ( .A(n24), .ZN(N16) );
  AOI22_X1 U64 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U65 ( .A(n25), .ZN(N17) );
  AOI22_X1 U66 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U67 ( .A(n21), .ZN(N13) );
  AOI22_X1 U68 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U69 ( .A(n29), .ZN(N20) );
  AOI22_X1 U70 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U71 ( .A(n30), .ZN(N21) );
  AOI22_X1 U72 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U73 ( .A(n20), .ZN(N12) );
  AOI22_X1 U74 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U75 ( .A(n19), .ZN(N11) );
  AOI22_X1 U76 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U77 ( .A(n18), .ZN(N10) );
  AOI22_X1 U78 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_58 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n5), .Z(n14) );
  BUF_X1 U4 ( .A(n4), .Z(n11) );
  BUF_X1 U5 ( .A(n4), .Z(n10) );
  BUF_X1 U6 ( .A(n6), .Z(n17) );
  BUF_X1 U7 ( .A(n4), .Z(n9) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n28), .ZN(N2) );
  INV_X1 U16 ( .A(n61), .ZN(N6) );
  AOI22_X1 U17 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U18 ( .A(n60), .ZN(N5) );
  AOI22_X1 U19 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U20 ( .A(n59), .ZN(N4) );
  AOI22_X1 U21 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U22 ( .A(n54), .ZN(N3) );
  AOI22_X1 U23 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U24 ( .A(n62), .ZN(N7) );
  AOI22_X1 U25 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U26 ( .A(n58), .ZN(N33) );
  AOI22_X1 U27 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U28 ( .A(n57), .ZN(N32) );
  AOI22_X1 U29 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U30 ( .A(n24), .ZN(N16) );
  AOI22_X1 U31 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U32 ( .A(n21), .ZN(N13) );
  AOI22_X1 U33 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U34 ( .A(n30), .ZN(N21) );
  AOI22_X1 U35 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U36 ( .A(n31), .ZN(N22) );
  AOI22_X1 U37 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U38 ( .A(n32), .ZN(N23) );
  AOI22_X1 U39 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U40 ( .A(n64), .ZN(N9) );
  AOI22_X1 U41 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U42 ( .A(n63), .ZN(N8) );
  AOI22_X1 U43 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U44 ( .A(n25), .ZN(N17) );
  AOI22_X1 U45 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U46 ( .A(n26), .ZN(N18) );
  AOI22_X1 U47 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U48 ( .A(n33), .ZN(N24) );
  AOI22_X1 U49 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U50 ( .A(n35), .ZN(N25) );
  AOI22_X1 U51 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U52 ( .A(n50), .ZN(N26) );
  AOI22_X1 U53 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U54 ( .A(n51), .ZN(N27) );
  AOI22_X1 U55 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U56 ( .A(n52), .ZN(N28) );
  AOI22_X1 U57 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U58 ( .A(n53), .ZN(N29) );
  AOI22_X1 U59 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U60 ( .A(n55), .ZN(N30) );
  AOI22_X1 U61 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U62 ( .A(n56), .ZN(N31) );
  AOI22_X1 U63 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U64 ( .A(n29), .ZN(N20) );
  AOI22_X1 U65 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U66 ( .A(n27), .ZN(N19) );
  AOI22_X1 U67 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U68 ( .A(n23), .ZN(N15) );
  AOI22_X1 U69 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U70 ( .A(n22), .ZN(N14) );
  AOI22_X1 U71 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U72 ( .A(n20), .ZN(N12) );
  AOI22_X1 U73 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U74 ( .A(n19), .ZN(N11) );
  AOI22_X1 U75 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U76 ( .A(n18), .ZN(N10) );
  AOI22_X1 U77 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U78 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_52 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n8) );
  INV_X1 U2 ( .A(n17), .ZN(n7) );
  AOI22_X1 U3 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U4 ( .A(n61), .ZN(N6) );
  INV_X1 U5 ( .A(n60), .ZN(N5) );
  INV_X1 U6 ( .A(n59), .ZN(N4) );
  INV_X1 U7 ( .A(n54), .ZN(N3) );
  INV_X1 U8 ( .A(n64), .ZN(N9) );
  INV_X1 U9 ( .A(n63), .ZN(N8) );
  INV_X1 U10 ( .A(n27), .ZN(N19) );
  INV_X1 U11 ( .A(n20), .ZN(N12) );
  INV_X1 U12 ( .A(n23), .ZN(N15) );
  INV_X1 U13 ( .A(n22), .ZN(N14) );
  INV_X1 U14 ( .A(n19), .ZN(N11) );
  INV_X1 U15 ( .A(n25), .ZN(N17) );
  INV_X1 U16 ( .A(n18), .ZN(N10) );
  INV_X1 U17 ( .A(n21), .ZN(N13) );
  INV_X1 U18 ( .A(n26), .ZN(N18) );
  BUF_X1 U19 ( .A(n4), .Z(n11) );
  BUF_X1 U20 ( .A(n5), .Z(n14) );
  BUF_X1 U21 ( .A(n6), .Z(n17) );
  INV_X1 U22 ( .A(n62), .ZN(N7) );
  INV_X1 U23 ( .A(n58), .ZN(N33) );
  INV_X1 U24 ( .A(n57), .ZN(N32) );
  INV_X1 U25 ( .A(n29), .ZN(N20) );
  INV_X1 U26 ( .A(n24), .ZN(N16) );
  INV_X1 U27 ( .A(n30), .ZN(N21) );
  INV_X1 U28 ( .A(n31), .ZN(N22) );
  INV_X1 U29 ( .A(n32), .ZN(N23) );
  INV_X1 U30 ( .A(n33), .ZN(N24) );
  INV_X1 U31 ( .A(n35), .ZN(N25) );
  INV_X1 U32 ( .A(n50), .ZN(N26) );
  INV_X1 U33 ( .A(n51), .ZN(N27) );
  INV_X1 U34 ( .A(n52), .ZN(N28) );
  INV_X1 U35 ( .A(n53), .ZN(N29) );
  INV_X1 U36 ( .A(n55), .ZN(N30) );
  INV_X1 U37 ( .A(n56), .ZN(N31) );
  BUF_X1 U38 ( .A(n4), .Z(n9) );
  BUF_X1 U39 ( .A(n6), .Z(n15) );
  BUF_X1 U40 ( .A(n4), .Z(n10) );
  BUF_X1 U41 ( .A(n6), .Z(n16) );
  BUF_X1 U42 ( .A(n5), .Z(n13) );
  BUF_X1 U43 ( .A(n5), .Z(n12) );
  AOI22_X1 U44 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U45 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U46 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U47 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U48 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U49 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U50 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U51 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U52 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U53 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U54 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U55 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U56 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U57 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U58 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U59 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U60 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U61 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U62 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  BUF_X1 U63 ( .A(sel), .Z(n6) );
  BUF_X1 U64 ( .A(sel), .Z(n5) );
  BUF_X1 U65 ( .A(sel), .Z(n4) );
  AOI22_X1 U66 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U67 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U68 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U69 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U70 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U71 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U72 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U73 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U74 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U75 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U77 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U78 ( .A(n28), .ZN(N2) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_48 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n59), .ZN(N4) );
  AOI22_X1 U16 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U17 ( .A(n60), .ZN(N5) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U19 ( .A(n61), .ZN(N6) );
  AOI22_X1 U20 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U21 ( .A(n62), .ZN(N7) );
  AOI22_X1 U22 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U23 ( .A(n63), .ZN(N8) );
  AOI22_X1 U24 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U25 ( .A(n64), .ZN(N9) );
  AOI22_X1 U26 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U31 ( .A(n28), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U33 ( .A(n54), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U35 ( .A(n18), .ZN(N10) );
  AOI22_X1 U36 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U37 ( .A(n19), .ZN(N11) );
  AOI22_X1 U38 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U39 ( .A(n20), .ZN(N12) );
  AOI22_X1 U40 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U41 ( .A(n21), .ZN(N13) );
  AOI22_X1 U42 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U43 ( .A(n22), .ZN(N14) );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U45 ( .A(n23), .ZN(N15) );
  AOI22_X1 U46 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U47 ( .A(n24), .ZN(N16) );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U49 ( .A(n25), .ZN(N17) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U51 ( .A(n26), .ZN(N18) );
  AOI22_X1 U52 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U53 ( .A(n27), .ZN(N19) );
  AOI22_X1 U54 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U55 ( .A(n29), .ZN(N20) );
  AOI22_X1 U56 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U57 ( .A(n30), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U59 ( .A(n31), .ZN(N22) );
  AOI22_X1 U60 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U61 ( .A(n32), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U63 ( .A(n33), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U65 ( .A(n35), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U67 ( .A(n50), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U69 ( .A(n51), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U71 ( .A(n52), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U73 ( .A(n53), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U75 ( .A(n55), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_47 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  AOI22_X1 U18 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U19 ( .A(n60), .ZN(N5) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U21 ( .A(n61), .ZN(N6) );
  AOI22_X1 U22 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U23 ( .A(n62), .ZN(N7) );
  AOI22_X1 U24 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U25 ( .A(n63), .ZN(N8) );
  AOI22_X1 U26 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U31 ( .A(n28), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U33 ( .A(n54), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U35 ( .A(n18), .ZN(N10) );
  AOI22_X1 U36 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U37 ( .A(n19), .ZN(N11) );
  AOI22_X1 U38 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U39 ( .A(n20), .ZN(N12) );
  AOI22_X1 U40 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U41 ( .A(n21), .ZN(N13) );
  AOI22_X1 U42 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U43 ( .A(n22), .ZN(N14) );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U45 ( .A(n23), .ZN(N15) );
  AOI22_X1 U46 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U47 ( .A(n24), .ZN(N16) );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U49 ( .A(n25), .ZN(N17) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U51 ( .A(n26), .ZN(N18) );
  AOI22_X1 U52 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U53 ( .A(n27), .ZN(N19) );
  AOI22_X1 U54 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U55 ( .A(n29), .ZN(N20) );
  AOI22_X1 U56 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U57 ( .A(n30), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U59 ( .A(n31), .ZN(N22) );
  AOI22_X1 U60 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U61 ( .A(n32), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U63 ( .A(n33), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U65 ( .A(n35), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U67 ( .A(n50), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U69 ( .A(n51), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U71 ( .A(n52), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U73 ( .A(n53), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U75 ( .A(n55), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_46 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  AOI22_X1 U18 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U19 ( .A(n60), .ZN(N5) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U21 ( .A(n61), .ZN(N6) );
  AOI22_X1 U22 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U23 ( .A(n62), .ZN(N7) );
  AOI22_X1 U24 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U25 ( .A(n63), .ZN(N8) );
  AOI22_X1 U26 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U31 ( .A(n28), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U33 ( .A(n54), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U35 ( .A(n18), .ZN(N10) );
  AOI22_X1 U36 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U37 ( .A(n19), .ZN(N11) );
  AOI22_X1 U38 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U39 ( .A(n20), .ZN(N12) );
  AOI22_X1 U40 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U41 ( .A(n21), .ZN(N13) );
  AOI22_X1 U42 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U43 ( .A(n22), .ZN(N14) );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U45 ( .A(n23), .ZN(N15) );
  AOI22_X1 U46 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U47 ( .A(n24), .ZN(N16) );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U49 ( .A(n25), .ZN(N17) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U51 ( .A(n26), .ZN(N18) );
  AOI22_X1 U52 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U53 ( .A(n27), .ZN(N19) );
  AOI22_X1 U54 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U55 ( .A(n29), .ZN(N20) );
  AOI22_X1 U56 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U57 ( .A(n30), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U59 ( .A(n31), .ZN(N22) );
  AOI22_X1 U60 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U61 ( .A(n32), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U63 ( .A(n33), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U65 ( .A(n35), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U67 ( .A(n50), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U69 ( .A(n51), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U71 ( .A(n52), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U73 ( .A(n53), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U75 ( .A(n55), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_45 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  AOI22_X1 U15 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U16 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U17 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U18 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U19 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U20 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U21 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U22 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U23 ( .A(n64), .ZN(N9) );
  AOI22_X1 U24 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U25 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U26 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U27 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U28 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U29 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U30 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U31 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U32 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U33 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U34 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U35 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U36 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U37 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U38 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U39 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U40 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U41 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U42 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U43 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U44 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U45 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U46 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U47 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U48 ( .A(n59), .ZN(N4) );
  INV_X1 U49 ( .A(n60), .ZN(N5) );
  INV_X1 U50 ( .A(n61), .ZN(N6) );
  INV_X1 U51 ( .A(n62), .ZN(N7) );
  INV_X1 U52 ( .A(n63), .ZN(N8) );
  INV_X1 U53 ( .A(n57), .ZN(N32) );
  INV_X1 U54 ( .A(n58), .ZN(N33) );
  INV_X1 U55 ( .A(n28), .ZN(N2) );
  INV_X1 U56 ( .A(n54), .ZN(N3) );
  INV_X1 U57 ( .A(n18), .ZN(N10) );
  INV_X1 U58 ( .A(n19), .ZN(N11) );
  INV_X1 U59 ( .A(n20), .ZN(N12) );
  INV_X1 U60 ( .A(n21), .ZN(N13) );
  INV_X1 U61 ( .A(n22), .ZN(N14) );
  INV_X1 U62 ( .A(n23), .ZN(N15) );
  INV_X1 U63 ( .A(n24), .ZN(N16) );
  INV_X1 U64 ( .A(n25), .ZN(N17) );
  INV_X1 U65 ( .A(n26), .ZN(N18) );
  INV_X1 U66 ( .A(n27), .ZN(N19) );
  INV_X1 U67 ( .A(n29), .ZN(N20) );
  INV_X1 U68 ( .A(n30), .ZN(N21) );
  INV_X1 U69 ( .A(n31), .ZN(N22) );
  INV_X1 U70 ( .A(n32), .ZN(N23) );
  INV_X1 U71 ( .A(n33), .ZN(N24) );
  INV_X1 U72 ( .A(n35), .ZN(N25) );
  INV_X1 U73 ( .A(n50), .ZN(N26) );
  INV_X1 U74 ( .A(n51), .ZN(N27) );
  INV_X1 U75 ( .A(n52), .ZN(N28) );
  INV_X1 U76 ( .A(n53), .ZN(N29) );
  INV_X1 U77 ( .A(n55), .ZN(N30) );
  INV_X1 U78 ( .A(n56), .ZN(N31) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_44 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n28), .ZN(N2) );
  AOI22_X1 U16 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U17 ( .A(n54), .ZN(N3) );
  AOI22_X1 U18 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U19 ( .A(n18), .ZN(N10) );
  AOI22_X1 U20 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U21 ( .A(n19), .ZN(N11) );
  AOI22_X1 U22 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U23 ( .A(n20), .ZN(N12) );
  AOI22_X1 U24 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U25 ( .A(n21), .ZN(N13) );
  AOI22_X1 U26 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U27 ( .A(n22), .ZN(N14) );
  AOI22_X1 U28 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U29 ( .A(n23), .ZN(N15) );
  AOI22_X1 U30 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U31 ( .A(n24), .ZN(N16) );
  AOI22_X1 U32 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U33 ( .A(n25), .ZN(N17) );
  AOI22_X1 U34 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U35 ( .A(n26), .ZN(N18) );
  AOI22_X1 U36 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U37 ( .A(n27), .ZN(N19) );
  AOI22_X1 U38 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U39 ( .A(n29), .ZN(N20) );
  AOI22_X1 U40 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U41 ( .A(n30), .ZN(N21) );
  AOI22_X1 U42 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U43 ( .A(n31), .ZN(N22) );
  AOI22_X1 U44 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U45 ( .A(n32), .ZN(N23) );
  AOI22_X1 U46 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U47 ( .A(n33), .ZN(N24) );
  AOI22_X1 U48 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U49 ( .A(n35), .ZN(N25) );
  AOI22_X1 U50 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U51 ( .A(n50), .ZN(N26) );
  AOI22_X1 U52 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U53 ( .A(n51), .ZN(N27) );
  AOI22_X1 U54 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U55 ( .A(n52), .ZN(N28) );
  AOI22_X1 U56 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U57 ( .A(n53), .ZN(N29) );
  AOI22_X1 U58 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U59 ( .A(n55), .ZN(N30) );
  AOI22_X1 U60 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U61 ( .A(n56), .ZN(N31) );
  AOI22_X1 U62 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U63 ( .A(n59), .ZN(N4) );
  AOI22_X1 U64 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U65 ( .A(n60), .ZN(N5) );
  AOI22_X1 U66 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U67 ( .A(n61), .ZN(N6) );
  AOI22_X1 U68 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U69 ( .A(n62), .ZN(N7) );
  AOI22_X1 U70 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U71 ( .A(n63), .ZN(N8) );
  AOI22_X1 U72 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U73 ( .A(n64), .ZN(N9) );
  AOI22_X1 U74 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U75 ( .A(n57), .ZN(N32) );
  AOI22_X1 U76 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U77 ( .A(n58), .ZN(N33) );
  AOI22_X1 U78 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_43 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  AOI22_X1 U18 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U19 ( .A(n60), .ZN(N5) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U21 ( .A(n61), .ZN(N6) );
  AOI22_X1 U22 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U23 ( .A(n62), .ZN(N7) );
  AOI22_X1 U24 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U25 ( .A(n63), .ZN(N8) );
  AOI22_X1 U26 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U31 ( .A(n28), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U33 ( .A(n54), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U35 ( .A(n18), .ZN(N10) );
  AOI22_X1 U36 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U37 ( .A(n19), .ZN(N11) );
  AOI22_X1 U38 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U39 ( .A(n20), .ZN(N12) );
  AOI22_X1 U40 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U41 ( .A(n21), .ZN(N13) );
  AOI22_X1 U42 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U43 ( .A(n22), .ZN(N14) );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U45 ( .A(n23), .ZN(N15) );
  AOI22_X1 U46 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U47 ( .A(n24), .ZN(N16) );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U49 ( .A(n25), .ZN(N17) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U51 ( .A(n26), .ZN(N18) );
  AOI22_X1 U52 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U53 ( .A(n27), .ZN(N19) );
  AOI22_X1 U54 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U55 ( .A(n29), .ZN(N20) );
  AOI22_X1 U56 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U57 ( .A(n30), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U59 ( .A(n31), .ZN(N22) );
  AOI22_X1 U60 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U61 ( .A(n32), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U63 ( .A(n33), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U65 ( .A(n35), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U67 ( .A(n50), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U69 ( .A(n51), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U71 ( .A(n52), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U73 ( .A(n53), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U75 ( .A(n55), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_42 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  AOI22_X1 U18 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U19 ( .A(n60), .ZN(N5) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U21 ( .A(n61), .ZN(N6) );
  AOI22_X1 U22 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U23 ( .A(n62), .ZN(N7) );
  AOI22_X1 U24 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U25 ( .A(n63), .ZN(N8) );
  AOI22_X1 U26 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U31 ( .A(n28), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U33 ( .A(n54), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U35 ( .A(n18), .ZN(N10) );
  AOI22_X1 U36 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U37 ( .A(n19), .ZN(N11) );
  AOI22_X1 U38 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U39 ( .A(n20), .ZN(N12) );
  AOI22_X1 U40 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U41 ( .A(n21), .ZN(N13) );
  AOI22_X1 U42 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U43 ( .A(n22), .ZN(N14) );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U45 ( .A(n23), .ZN(N15) );
  AOI22_X1 U46 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U47 ( .A(n24), .ZN(N16) );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U49 ( .A(n25), .ZN(N17) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U51 ( .A(n26), .ZN(N18) );
  AOI22_X1 U52 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U53 ( .A(n27), .ZN(N19) );
  AOI22_X1 U54 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U55 ( .A(n29), .ZN(N20) );
  AOI22_X1 U56 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U57 ( .A(n30), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U59 ( .A(n31), .ZN(N22) );
  AOI22_X1 U60 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U61 ( .A(n32), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U63 ( .A(n33), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U65 ( .A(n35), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U67 ( .A(n50), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U69 ( .A(n51), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U71 ( .A(n52), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U73 ( .A(n53), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U75 ( .A(n55), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_41 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  AOI22_X1 U15 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U16 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U17 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U18 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U19 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U20 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U21 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U22 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U23 ( .A(n64), .ZN(N9) );
  AOI22_X1 U24 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U25 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U26 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U27 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U28 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U29 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U30 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U31 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U32 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U33 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U34 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U35 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U36 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U37 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U38 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U39 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U40 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U41 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U42 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U43 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U44 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U45 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U46 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U47 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U48 ( .A(n59), .ZN(N4) );
  INV_X1 U49 ( .A(n60), .ZN(N5) );
  INV_X1 U50 ( .A(n61), .ZN(N6) );
  INV_X1 U51 ( .A(n62), .ZN(N7) );
  INV_X1 U52 ( .A(n63), .ZN(N8) );
  INV_X1 U53 ( .A(n57), .ZN(N32) );
  INV_X1 U54 ( .A(n58), .ZN(N33) );
  INV_X1 U55 ( .A(n28), .ZN(N2) );
  INV_X1 U56 ( .A(n54), .ZN(N3) );
  INV_X1 U57 ( .A(n18), .ZN(N10) );
  INV_X1 U58 ( .A(n19), .ZN(N11) );
  INV_X1 U59 ( .A(n20), .ZN(N12) );
  INV_X1 U60 ( .A(n21), .ZN(N13) );
  INV_X1 U61 ( .A(n22), .ZN(N14) );
  INV_X1 U62 ( .A(n23), .ZN(N15) );
  INV_X1 U63 ( .A(n24), .ZN(N16) );
  INV_X1 U64 ( .A(n25), .ZN(N17) );
  INV_X1 U65 ( .A(n26), .ZN(N18) );
  INV_X1 U66 ( .A(n27), .ZN(N19) );
  INV_X1 U67 ( .A(n29), .ZN(N20) );
  INV_X1 U68 ( .A(n30), .ZN(N21) );
  INV_X1 U69 ( .A(n31), .ZN(N22) );
  INV_X1 U70 ( .A(n32), .ZN(N23) );
  INV_X1 U71 ( .A(n33), .ZN(N24) );
  INV_X1 U72 ( .A(n35), .ZN(N25) );
  INV_X1 U73 ( .A(n50), .ZN(N26) );
  INV_X1 U74 ( .A(n51), .ZN(N27) );
  INV_X1 U75 ( .A(n52), .ZN(N28) );
  INV_X1 U76 ( .A(n53), .ZN(N29) );
  INV_X1 U77 ( .A(n55), .ZN(N30) );
  INV_X1 U78 ( .A(n56), .ZN(N31) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_40 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n28), .ZN(N2) );
  AOI22_X1 U16 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U17 ( .A(n54), .ZN(N3) );
  AOI22_X1 U18 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U19 ( .A(n18), .ZN(N10) );
  AOI22_X1 U20 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U21 ( .A(n19), .ZN(N11) );
  AOI22_X1 U22 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U23 ( .A(n20), .ZN(N12) );
  AOI22_X1 U24 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U25 ( .A(n21), .ZN(N13) );
  AOI22_X1 U26 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U27 ( .A(n22), .ZN(N14) );
  AOI22_X1 U28 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U29 ( .A(n23), .ZN(N15) );
  AOI22_X1 U30 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U31 ( .A(n24), .ZN(N16) );
  AOI22_X1 U32 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U33 ( .A(n25), .ZN(N17) );
  AOI22_X1 U34 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U35 ( .A(n26), .ZN(N18) );
  AOI22_X1 U36 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U37 ( .A(n27), .ZN(N19) );
  AOI22_X1 U38 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U39 ( .A(n29), .ZN(N20) );
  AOI22_X1 U40 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U41 ( .A(n30), .ZN(N21) );
  AOI22_X1 U42 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U43 ( .A(n31), .ZN(N22) );
  AOI22_X1 U44 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U45 ( .A(n32), .ZN(N23) );
  AOI22_X1 U46 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U47 ( .A(n33), .ZN(N24) );
  AOI22_X1 U48 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U49 ( .A(n35), .ZN(N25) );
  AOI22_X1 U50 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U51 ( .A(n50), .ZN(N26) );
  AOI22_X1 U52 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U53 ( .A(n51), .ZN(N27) );
  AOI22_X1 U54 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U55 ( .A(n52), .ZN(N28) );
  AOI22_X1 U56 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U57 ( .A(n53), .ZN(N29) );
  AOI22_X1 U58 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U59 ( .A(n55), .ZN(N30) );
  AOI22_X1 U60 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U61 ( .A(n56), .ZN(N31) );
  AOI22_X1 U62 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U63 ( .A(n59), .ZN(N4) );
  AOI22_X1 U64 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U65 ( .A(n60), .ZN(N5) );
  AOI22_X1 U66 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U67 ( .A(n61), .ZN(N6) );
  AOI22_X1 U68 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U69 ( .A(n62), .ZN(N7) );
  AOI22_X1 U70 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U71 ( .A(n63), .ZN(N8) );
  AOI22_X1 U72 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U73 ( .A(n64), .ZN(N9) );
  AOI22_X1 U74 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U75 ( .A(n57), .ZN(N32) );
  AOI22_X1 U76 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U77 ( .A(n58), .ZN(N33) );
  AOI22_X1 U78 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_39 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  AOI22_X1 U18 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U19 ( .A(n60), .ZN(N5) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U21 ( .A(n61), .ZN(N6) );
  AOI22_X1 U22 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U23 ( .A(n62), .ZN(N7) );
  AOI22_X1 U24 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U25 ( .A(n63), .ZN(N8) );
  AOI22_X1 U26 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U31 ( .A(n28), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U33 ( .A(n54), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U35 ( .A(n18), .ZN(N10) );
  AOI22_X1 U36 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U37 ( .A(n19), .ZN(N11) );
  AOI22_X1 U38 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U39 ( .A(n20), .ZN(N12) );
  AOI22_X1 U40 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U41 ( .A(n21), .ZN(N13) );
  AOI22_X1 U42 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U43 ( .A(n22), .ZN(N14) );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U45 ( .A(n23), .ZN(N15) );
  AOI22_X1 U46 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U47 ( .A(n24), .ZN(N16) );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U49 ( .A(n25), .ZN(N17) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U51 ( .A(n26), .ZN(N18) );
  AOI22_X1 U52 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U53 ( .A(n27), .ZN(N19) );
  AOI22_X1 U54 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U55 ( .A(n29), .ZN(N20) );
  AOI22_X1 U56 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U57 ( .A(n30), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U59 ( .A(n31), .ZN(N22) );
  AOI22_X1 U60 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U61 ( .A(n32), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U63 ( .A(n33), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U65 ( .A(n35), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U67 ( .A(n50), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U69 ( .A(n51), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U71 ( .A(n52), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U73 ( .A(n53), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U75 ( .A(n55), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_38 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  AOI22_X1 U18 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U19 ( .A(n60), .ZN(N5) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U21 ( .A(n61), .ZN(N6) );
  AOI22_X1 U22 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U23 ( .A(n62), .ZN(N7) );
  AOI22_X1 U24 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U25 ( .A(n63), .ZN(N8) );
  AOI22_X1 U26 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U31 ( .A(n28), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U33 ( .A(n54), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U35 ( .A(n18), .ZN(N10) );
  AOI22_X1 U36 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U37 ( .A(n19), .ZN(N11) );
  AOI22_X1 U38 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U39 ( .A(n20), .ZN(N12) );
  AOI22_X1 U40 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U41 ( .A(n21), .ZN(N13) );
  AOI22_X1 U42 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U43 ( .A(n22), .ZN(N14) );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U45 ( .A(n23), .ZN(N15) );
  AOI22_X1 U46 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U47 ( .A(n24), .ZN(N16) );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U49 ( .A(n25), .ZN(N17) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U51 ( .A(n26), .ZN(N18) );
  AOI22_X1 U52 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U53 ( .A(n27), .ZN(N19) );
  AOI22_X1 U54 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U55 ( .A(n29), .ZN(N20) );
  AOI22_X1 U56 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U57 ( .A(n30), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U59 ( .A(n31), .ZN(N22) );
  AOI22_X1 U60 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U61 ( .A(n32), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U63 ( .A(n33), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U65 ( .A(n35), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U67 ( .A(n50), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U69 ( .A(n51), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U71 ( .A(n52), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U73 ( .A(n53), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U75 ( .A(n55), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_37 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  AOI22_X1 U15 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U16 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U17 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U18 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U19 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U20 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U21 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U22 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U23 ( .A(n64), .ZN(N9) );
  AOI22_X1 U24 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U25 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U26 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U27 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U28 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U29 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U30 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U31 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U32 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U33 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U34 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U35 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U36 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U37 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U38 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U39 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U40 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U41 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U42 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U43 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U44 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U45 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U46 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U47 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U48 ( .A(n59), .ZN(N4) );
  INV_X1 U49 ( .A(n60), .ZN(N5) );
  INV_X1 U50 ( .A(n61), .ZN(N6) );
  INV_X1 U51 ( .A(n62), .ZN(N7) );
  INV_X1 U52 ( .A(n63), .ZN(N8) );
  INV_X1 U53 ( .A(n57), .ZN(N32) );
  INV_X1 U54 ( .A(n58), .ZN(N33) );
  INV_X1 U55 ( .A(n28), .ZN(N2) );
  INV_X1 U56 ( .A(n54), .ZN(N3) );
  INV_X1 U57 ( .A(n18), .ZN(N10) );
  INV_X1 U58 ( .A(n19), .ZN(N11) );
  INV_X1 U59 ( .A(n20), .ZN(N12) );
  INV_X1 U60 ( .A(n21), .ZN(N13) );
  INV_X1 U61 ( .A(n22), .ZN(N14) );
  INV_X1 U62 ( .A(n23), .ZN(N15) );
  INV_X1 U63 ( .A(n24), .ZN(N16) );
  INV_X1 U64 ( .A(n25), .ZN(N17) );
  INV_X1 U65 ( .A(n26), .ZN(N18) );
  INV_X1 U66 ( .A(n27), .ZN(N19) );
  INV_X1 U67 ( .A(n29), .ZN(N20) );
  INV_X1 U68 ( .A(n30), .ZN(N21) );
  INV_X1 U69 ( .A(n31), .ZN(N22) );
  INV_X1 U70 ( .A(n32), .ZN(N23) );
  INV_X1 U71 ( .A(n33), .ZN(N24) );
  INV_X1 U72 ( .A(n35), .ZN(N25) );
  INV_X1 U73 ( .A(n50), .ZN(N26) );
  INV_X1 U74 ( .A(n51), .ZN(N27) );
  INV_X1 U75 ( .A(n52), .ZN(N28) );
  INV_X1 U76 ( .A(n53), .ZN(N29) );
  INV_X1 U77 ( .A(n55), .ZN(N30) );
  INV_X1 U78 ( .A(n56), .ZN(N31) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_36 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U17 ( .A(n28), .ZN(N2) );
  AOI22_X1 U18 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U19 ( .A(n54), .ZN(N3) );
  AOI22_X1 U20 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U21 ( .A(n18), .ZN(N10) );
  AOI22_X1 U22 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U23 ( .A(n19), .ZN(N11) );
  AOI22_X1 U24 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U25 ( .A(n20), .ZN(N12) );
  AOI22_X1 U26 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U27 ( .A(n21), .ZN(N13) );
  AOI22_X1 U28 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U29 ( .A(n22), .ZN(N14) );
  AOI22_X1 U30 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U31 ( .A(n23), .ZN(N15) );
  AOI22_X1 U32 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U33 ( .A(n24), .ZN(N16) );
  AOI22_X1 U34 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U35 ( .A(n25), .ZN(N17) );
  AOI22_X1 U36 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U37 ( .A(n26), .ZN(N18) );
  AOI22_X1 U38 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U39 ( .A(n27), .ZN(N19) );
  AOI22_X1 U40 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U41 ( .A(n29), .ZN(N20) );
  AOI22_X1 U42 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U43 ( .A(n30), .ZN(N21) );
  AOI22_X1 U44 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U45 ( .A(n31), .ZN(N22) );
  AOI22_X1 U46 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U47 ( .A(n32), .ZN(N23) );
  AOI22_X1 U48 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U49 ( .A(n33), .ZN(N24) );
  AOI22_X1 U50 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U51 ( .A(n35), .ZN(N25) );
  AOI22_X1 U52 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U53 ( .A(n50), .ZN(N26) );
  AOI22_X1 U54 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U55 ( .A(n51), .ZN(N27) );
  AOI22_X1 U56 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U57 ( .A(n52), .ZN(N28) );
  AOI22_X1 U58 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U59 ( .A(n53), .ZN(N29) );
  AOI22_X1 U60 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U61 ( .A(n55), .ZN(N30) );
  AOI22_X1 U62 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U63 ( .A(n56), .ZN(N31) );
  AOI22_X1 U64 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U65 ( .A(n59), .ZN(N4) );
  AOI22_X1 U66 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U67 ( .A(n60), .ZN(N5) );
  AOI22_X1 U68 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U69 ( .A(n61), .ZN(N6) );
  AOI22_X1 U70 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U71 ( .A(n62), .ZN(N7) );
  AOI22_X1 U72 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U73 ( .A(n63), .ZN(N8) );
  AOI22_X1 U74 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U75 ( .A(n57), .ZN(N32) );
  AOI22_X1 U76 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U77 ( .A(n58), .ZN(N33) );
  AOI22_X1 U78 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_35 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  AOI22_X1 U18 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U19 ( .A(n60), .ZN(N5) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U21 ( .A(n61), .ZN(N6) );
  AOI22_X1 U22 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U23 ( .A(n62), .ZN(N7) );
  AOI22_X1 U24 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U25 ( .A(n63), .ZN(N8) );
  AOI22_X1 U26 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U31 ( .A(n28), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U33 ( .A(n54), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U35 ( .A(n18), .ZN(N10) );
  AOI22_X1 U36 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U37 ( .A(n19), .ZN(N11) );
  AOI22_X1 U38 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U39 ( .A(n20), .ZN(N12) );
  AOI22_X1 U40 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U41 ( .A(n21), .ZN(N13) );
  AOI22_X1 U42 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U43 ( .A(n22), .ZN(N14) );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U45 ( .A(n23), .ZN(N15) );
  AOI22_X1 U46 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U47 ( .A(n24), .ZN(N16) );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U49 ( .A(n25), .ZN(N17) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U51 ( .A(n26), .ZN(N18) );
  AOI22_X1 U52 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U53 ( .A(n27), .ZN(N19) );
  AOI22_X1 U54 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U55 ( .A(n29), .ZN(N20) );
  AOI22_X1 U56 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U57 ( .A(n30), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U59 ( .A(n31), .ZN(N22) );
  AOI22_X1 U60 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U61 ( .A(n32), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U63 ( .A(n33), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U65 ( .A(n35), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U67 ( .A(n50), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U69 ( .A(n51), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U71 ( .A(n52), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U73 ( .A(n53), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U75 ( .A(n55), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_34 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  AOI22_X1 U18 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U19 ( .A(n60), .ZN(N5) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U21 ( .A(n61), .ZN(N6) );
  AOI22_X1 U22 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U23 ( .A(n62), .ZN(N7) );
  AOI22_X1 U24 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U25 ( .A(n63), .ZN(N8) );
  AOI22_X1 U26 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U31 ( .A(n28), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U33 ( .A(n54), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U35 ( .A(n18), .ZN(N10) );
  AOI22_X1 U36 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U37 ( .A(n19), .ZN(N11) );
  AOI22_X1 U38 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U39 ( .A(n20), .ZN(N12) );
  AOI22_X1 U40 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U41 ( .A(n21), .ZN(N13) );
  AOI22_X1 U42 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U43 ( .A(n22), .ZN(N14) );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U45 ( .A(n23), .ZN(N15) );
  AOI22_X1 U46 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U47 ( .A(n24), .ZN(N16) );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U49 ( .A(n25), .ZN(N17) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U51 ( .A(n26), .ZN(N18) );
  AOI22_X1 U52 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U53 ( .A(n27), .ZN(N19) );
  AOI22_X1 U54 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U55 ( .A(n29), .ZN(N20) );
  AOI22_X1 U56 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U57 ( .A(n30), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U59 ( .A(n31), .ZN(N22) );
  AOI22_X1 U60 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U61 ( .A(n32), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U63 ( .A(n33), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U65 ( .A(n35), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U67 ( .A(n50), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U69 ( .A(n51), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U71 ( .A(n52), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U73 ( .A(n53), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U75 ( .A(n55), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_33 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  AOI22_X1 U15 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U16 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U17 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U18 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U19 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U20 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U21 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U22 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U23 ( .A(n64), .ZN(N9) );
  AOI22_X1 U24 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U25 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U26 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U27 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U28 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U29 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U30 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U31 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U32 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U33 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U34 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U35 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U36 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U37 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U38 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U39 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U40 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U41 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U42 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U43 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U44 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U45 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U46 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U47 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U48 ( .A(n59), .ZN(N4) );
  INV_X1 U49 ( .A(n60), .ZN(N5) );
  INV_X1 U50 ( .A(n61), .ZN(N6) );
  INV_X1 U51 ( .A(n62), .ZN(N7) );
  INV_X1 U52 ( .A(n63), .ZN(N8) );
  INV_X1 U53 ( .A(n57), .ZN(N32) );
  INV_X1 U54 ( .A(n58), .ZN(N33) );
  INV_X1 U55 ( .A(n28), .ZN(N2) );
  INV_X1 U56 ( .A(n54), .ZN(N3) );
  INV_X1 U57 ( .A(n18), .ZN(N10) );
  INV_X1 U58 ( .A(n19), .ZN(N11) );
  INV_X1 U59 ( .A(n20), .ZN(N12) );
  INV_X1 U60 ( .A(n21), .ZN(N13) );
  INV_X1 U61 ( .A(n22), .ZN(N14) );
  INV_X1 U62 ( .A(n23), .ZN(N15) );
  INV_X1 U63 ( .A(n24), .ZN(N16) );
  INV_X1 U64 ( .A(n25), .ZN(N17) );
  INV_X1 U65 ( .A(n26), .ZN(N18) );
  INV_X1 U66 ( .A(n27), .ZN(N19) );
  INV_X1 U67 ( .A(n29), .ZN(N20) );
  INV_X1 U68 ( .A(n30), .ZN(N21) );
  INV_X1 U69 ( .A(n31), .ZN(N22) );
  INV_X1 U70 ( .A(n32), .ZN(N23) );
  INV_X1 U71 ( .A(n33), .ZN(N24) );
  INV_X1 U72 ( .A(n35), .ZN(N25) );
  INV_X1 U73 ( .A(n50), .ZN(N26) );
  INV_X1 U74 ( .A(n51), .ZN(N27) );
  INV_X1 U75 ( .A(n52), .ZN(N28) );
  INV_X1 U76 ( .A(n53), .ZN(N29) );
  INV_X1 U77 ( .A(n55), .ZN(N30) );
  INV_X1 U78 ( .A(n56), .ZN(N31) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_32 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n6), .Z(n17) );
  BUF_X1 U4 ( .A(n4), .Z(n9) );
  BUF_X1 U5 ( .A(n6), .Z(n15) );
  BUF_X1 U6 ( .A(n5), .Z(n14) );
  BUF_X1 U7 ( .A(n5), .Z(n12) );
  BUF_X1 U8 ( .A(n4), .Z(n11) );
  BUF_X1 U9 ( .A(n5), .Z(n13) );
  BUF_X1 U10 ( .A(n4), .Z(n10) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  AOI22_X1 U18 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U19 ( .A(n60), .ZN(N5) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U21 ( .A(n61), .ZN(N6) );
  AOI22_X1 U22 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U23 ( .A(n62), .ZN(N7) );
  AOI22_X1 U24 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U25 ( .A(n63), .ZN(N8) );
  AOI22_X1 U26 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U31 ( .A(n28), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U33 ( .A(n54), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U35 ( .A(n21), .ZN(N13) );
  AOI22_X1 U36 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U37 ( .A(n22), .ZN(N14) );
  AOI22_X1 U38 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U39 ( .A(n23), .ZN(N15) );
  AOI22_X1 U40 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U41 ( .A(n24), .ZN(N16) );
  AOI22_X1 U42 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U43 ( .A(n25), .ZN(N17) );
  AOI22_X1 U44 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U45 ( .A(n26), .ZN(N18) );
  AOI22_X1 U46 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U47 ( .A(n27), .ZN(N19) );
  AOI22_X1 U48 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U49 ( .A(n29), .ZN(N20) );
  AOI22_X1 U50 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U51 ( .A(n30), .ZN(N21) );
  AOI22_X1 U52 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U53 ( .A(n31), .ZN(N22) );
  AOI22_X1 U54 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U55 ( .A(n32), .ZN(N23) );
  AOI22_X1 U56 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U57 ( .A(n33), .ZN(N24) );
  AOI22_X1 U58 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U59 ( .A(n35), .ZN(N25) );
  AOI22_X1 U60 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U61 ( .A(n50), .ZN(N26) );
  AOI22_X1 U62 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U63 ( .A(n51), .ZN(N27) );
  AOI22_X1 U64 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U65 ( .A(n52), .ZN(N28) );
  AOI22_X1 U66 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U67 ( .A(n53), .ZN(N29) );
  AOI22_X1 U68 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U69 ( .A(n55), .ZN(N30) );
  AOI22_X1 U70 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U71 ( .A(n56), .ZN(N31) );
  AOI22_X1 U72 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U73 ( .A(n18), .ZN(N10) );
  AOI22_X1 U74 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U75 ( .A(n19), .ZN(N11) );
  AOI22_X1 U76 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U77 ( .A(n20), .ZN(N12) );
  AOI22_X1 U78 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_31 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n6), .Z(n17) );
  BUF_X1 U4 ( .A(n4), .Z(n9) );
  BUF_X1 U5 ( .A(n6), .Z(n15) );
  BUF_X1 U6 ( .A(n5), .Z(n14) );
  BUF_X1 U7 ( .A(n5), .Z(n12) );
  BUF_X1 U8 ( .A(n4), .Z(n11) );
  BUF_X1 U9 ( .A(n5), .Z(n13) );
  BUF_X1 U10 ( .A(n4), .Z(n10) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  INV_X1 U16 ( .A(n59), .ZN(N4) );
  INV_X1 U17 ( .A(n60), .ZN(N5) );
  INV_X1 U18 ( .A(n61), .ZN(N6) );
  INV_X1 U19 ( .A(n62), .ZN(N7) );
  INV_X1 U20 ( .A(n63), .ZN(N8) );
  INV_X1 U21 ( .A(n57), .ZN(N32) );
  INV_X1 U22 ( .A(n58), .ZN(N33) );
  INV_X1 U23 ( .A(n28), .ZN(N2) );
  INV_X1 U24 ( .A(n54), .ZN(N3) );
  INV_X1 U25 ( .A(n21), .ZN(N13) );
  INV_X1 U26 ( .A(n22), .ZN(N14) );
  INV_X1 U27 ( .A(n23), .ZN(N15) );
  INV_X1 U28 ( .A(n24), .ZN(N16) );
  INV_X1 U29 ( .A(n25), .ZN(N17) );
  INV_X1 U30 ( .A(n26), .ZN(N18) );
  INV_X1 U31 ( .A(n27), .ZN(N19) );
  INV_X1 U32 ( .A(n29), .ZN(N20) );
  INV_X1 U33 ( .A(n30), .ZN(N21) );
  INV_X1 U34 ( .A(n31), .ZN(N22) );
  INV_X1 U35 ( .A(n32), .ZN(N23) );
  INV_X1 U36 ( .A(n33), .ZN(N24) );
  INV_X1 U37 ( .A(n35), .ZN(N25) );
  INV_X1 U38 ( .A(n50), .ZN(N26) );
  INV_X1 U39 ( .A(n51), .ZN(N27) );
  INV_X1 U40 ( .A(n52), .ZN(N28) );
  INV_X1 U41 ( .A(n53), .ZN(N29) );
  INV_X1 U42 ( .A(n55), .ZN(N30) );
  INV_X1 U43 ( .A(n56), .ZN(N31) );
  INV_X1 U44 ( .A(n18), .ZN(N10) );
  INV_X1 U45 ( .A(n19), .ZN(N11) );
  INV_X1 U46 ( .A(n20), .ZN(N12) );
  AOI22_X1 U47 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U48 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U49 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U50 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U51 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U52 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U53 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U54 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U55 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U56 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U57 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U58 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U59 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U60 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U61 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U62 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U63 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U64 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U65 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U66 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_30 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n6), .Z(n17) );
  BUF_X1 U4 ( .A(n4), .Z(n9) );
  BUF_X1 U5 ( .A(n6), .Z(n15) );
  BUF_X1 U6 ( .A(n5), .Z(n14) );
  BUF_X1 U7 ( .A(n5), .Z(n12) );
  BUF_X1 U8 ( .A(n4), .Z(n11) );
  BUF_X1 U9 ( .A(n5), .Z(n13) );
  BUF_X1 U10 ( .A(n4), .Z(n10) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  AOI22_X1 U18 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U19 ( .A(n60), .ZN(N5) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U21 ( .A(n61), .ZN(N6) );
  AOI22_X1 U22 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U23 ( .A(n62), .ZN(N7) );
  AOI22_X1 U24 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U25 ( .A(n63), .ZN(N8) );
  AOI22_X1 U26 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U31 ( .A(n28), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U33 ( .A(n54), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U35 ( .A(n21), .ZN(N13) );
  AOI22_X1 U36 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U37 ( .A(n22), .ZN(N14) );
  AOI22_X1 U38 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U39 ( .A(n23), .ZN(N15) );
  AOI22_X1 U40 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U41 ( .A(n24), .ZN(N16) );
  AOI22_X1 U42 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U43 ( .A(n25), .ZN(N17) );
  AOI22_X1 U44 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U45 ( .A(n26), .ZN(N18) );
  AOI22_X1 U46 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U47 ( .A(n27), .ZN(N19) );
  AOI22_X1 U48 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U49 ( .A(n29), .ZN(N20) );
  AOI22_X1 U50 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U51 ( .A(n30), .ZN(N21) );
  AOI22_X1 U52 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U53 ( .A(n31), .ZN(N22) );
  AOI22_X1 U54 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U55 ( .A(n32), .ZN(N23) );
  AOI22_X1 U56 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U57 ( .A(n33), .ZN(N24) );
  AOI22_X1 U58 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U59 ( .A(n35), .ZN(N25) );
  AOI22_X1 U60 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U61 ( .A(n50), .ZN(N26) );
  AOI22_X1 U62 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U63 ( .A(n51), .ZN(N27) );
  AOI22_X1 U64 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U65 ( .A(n52), .ZN(N28) );
  AOI22_X1 U66 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U67 ( .A(n53), .ZN(N29) );
  AOI22_X1 U68 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U69 ( .A(n55), .ZN(N30) );
  AOI22_X1 U70 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U71 ( .A(n56), .ZN(N31) );
  AOI22_X1 U72 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U73 ( .A(n18), .ZN(N10) );
  AOI22_X1 U74 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U75 ( .A(n19), .ZN(N11) );
  AOI22_X1 U76 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U77 ( .A(n20), .ZN(N12) );
  AOI22_X1 U78 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_29 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n6), .Z(n17) );
  BUF_X1 U4 ( .A(n4), .Z(n9) );
  BUF_X1 U5 ( .A(n6), .Z(n15) );
  BUF_X1 U6 ( .A(n5), .Z(n14) );
  BUF_X1 U7 ( .A(n5), .Z(n12) );
  BUF_X1 U8 ( .A(n4), .Z(n11) );
  BUF_X1 U9 ( .A(n5), .Z(n13) );
  BUF_X1 U10 ( .A(n4), .Z(n10) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  INV_X1 U16 ( .A(n59), .ZN(N4) );
  INV_X1 U17 ( .A(n60), .ZN(N5) );
  INV_X1 U18 ( .A(n61), .ZN(N6) );
  INV_X1 U19 ( .A(n62), .ZN(N7) );
  INV_X1 U20 ( .A(n63), .ZN(N8) );
  INV_X1 U21 ( .A(n57), .ZN(N32) );
  INV_X1 U22 ( .A(n58), .ZN(N33) );
  INV_X1 U23 ( .A(n28), .ZN(N2) );
  INV_X1 U24 ( .A(n54), .ZN(N3) );
  INV_X1 U25 ( .A(n21), .ZN(N13) );
  INV_X1 U26 ( .A(n22), .ZN(N14) );
  INV_X1 U27 ( .A(n23), .ZN(N15) );
  INV_X1 U28 ( .A(n24), .ZN(N16) );
  INV_X1 U29 ( .A(n25), .ZN(N17) );
  INV_X1 U30 ( .A(n26), .ZN(N18) );
  INV_X1 U31 ( .A(n27), .ZN(N19) );
  INV_X1 U32 ( .A(n29), .ZN(N20) );
  INV_X1 U33 ( .A(n30), .ZN(N21) );
  INV_X1 U34 ( .A(n31), .ZN(N22) );
  INV_X1 U35 ( .A(n32), .ZN(N23) );
  INV_X1 U36 ( .A(n33), .ZN(N24) );
  INV_X1 U37 ( .A(n35), .ZN(N25) );
  INV_X1 U38 ( .A(n50), .ZN(N26) );
  INV_X1 U39 ( .A(n51), .ZN(N27) );
  INV_X1 U40 ( .A(n52), .ZN(N28) );
  INV_X1 U41 ( .A(n53), .ZN(N29) );
  INV_X1 U42 ( .A(n55), .ZN(N30) );
  INV_X1 U43 ( .A(n56), .ZN(N31) );
  INV_X1 U44 ( .A(n18), .ZN(N10) );
  INV_X1 U45 ( .A(n19), .ZN(N11) );
  INV_X1 U46 ( .A(n20), .ZN(N12) );
  AOI22_X1 U47 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U48 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U49 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U50 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U51 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U52 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U53 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U54 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U55 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U56 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U57 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U58 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U59 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U60 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U61 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U62 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U63 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U64 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U65 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U66 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_28 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n6), .Z(n17) );
  BUF_X1 U4 ( .A(n4), .Z(n9) );
  BUF_X1 U5 ( .A(n6), .Z(n15) );
  BUF_X1 U6 ( .A(n5), .Z(n14) );
  BUF_X1 U7 ( .A(n5), .Z(n12) );
  BUF_X1 U8 ( .A(n4), .Z(n11) );
  BUF_X1 U9 ( .A(n5), .Z(n13) );
  BUF_X1 U10 ( .A(n4), .Z(n10) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  AOI22_X1 U18 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U19 ( .A(n60), .ZN(N5) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U21 ( .A(n61), .ZN(N6) );
  AOI22_X1 U22 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U23 ( .A(n62), .ZN(N7) );
  AOI22_X1 U24 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U25 ( .A(n63), .ZN(N8) );
  AOI22_X1 U26 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U31 ( .A(n28), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U33 ( .A(n54), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U35 ( .A(n21), .ZN(N13) );
  AOI22_X1 U36 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U37 ( .A(n22), .ZN(N14) );
  AOI22_X1 U38 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U39 ( .A(n23), .ZN(N15) );
  AOI22_X1 U40 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U41 ( .A(n24), .ZN(N16) );
  AOI22_X1 U42 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U43 ( .A(n25), .ZN(N17) );
  AOI22_X1 U44 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U45 ( .A(n26), .ZN(N18) );
  AOI22_X1 U46 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U47 ( .A(n27), .ZN(N19) );
  AOI22_X1 U48 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U49 ( .A(n29), .ZN(N20) );
  AOI22_X1 U50 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U51 ( .A(n30), .ZN(N21) );
  AOI22_X1 U52 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U53 ( .A(n31), .ZN(N22) );
  AOI22_X1 U54 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U55 ( .A(n32), .ZN(N23) );
  AOI22_X1 U56 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U57 ( .A(n33), .ZN(N24) );
  AOI22_X1 U58 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U59 ( .A(n35), .ZN(N25) );
  AOI22_X1 U60 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U61 ( .A(n50), .ZN(N26) );
  AOI22_X1 U62 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U63 ( .A(n51), .ZN(N27) );
  AOI22_X1 U64 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U65 ( .A(n52), .ZN(N28) );
  AOI22_X1 U66 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U67 ( .A(n53), .ZN(N29) );
  AOI22_X1 U68 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U69 ( .A(n55), .ZN(N30) );
  AOI22_X1 U70 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U71 ( .A(n56), .ZN(N31) );
  AOI22_X1 U72 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U73 ( .A(n18), .ZN(N10) );
  AOI22_X1 U74 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U75 ( .A(n19), .ZN(N11) );
  AOI22_X1 U76 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U77 ( .A(n20), .ZN(N12) );
  AOI22_X1 U78 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_27 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n6), .Z(n17) );
  BUF_X1 U4 ( .A(n4), .Z(n9) );
  BUF_X1 U5 ( .A(n6), .Z(n15) );
  BUF_X1 U6 ( .A(n5), .Z(n14) );
  BUF_X1 U7 ( .A(n5), .Z(n12) );
  BUF_X1 U8 ( .A(n4), .Z(n11) );
  BUF_X1 U9 ( .A(n5), .Z(n13) );
  BUF_X1 U10 ( .A(n4), .Z(n10) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  INV_X1 U16 ( .A(n59), .ZN(N4) );
  INV_X1 U17 ( .A(n60), .ZN(N5) );
  INV_X1 U18 ( .A(n61), .ZN(N6) );
  INV_X1 U19 ( .A(n62), .ZN(N7) );
  INV_X1 U20 ( .A(n63), .ZN(N8) );
  INV_X1 U21 ( .A(n57), .ZN(N32) );
  INV_X1 U22 ( .A(n58), .ZN(N33) );
  INV_X1 U23 ( .A(n28), .ZN(N2) );
  INV_X1 U24 ( .A(n54), .ZN(N3) );
  INV_X1 U25 ( .A(n21), .ZN(N13) );
  INV_X1 U26 ( .A(n22), .ZN(N14) );
  INV_X1 U27 ( .A(n23), .ZN(N15) );
  INV_X1 U28 ( .A(n24), .ZN(N16) );
  INV_X1 U29 ( .A(n25), .ZN(N17) );
  INV_X1 U30 ( .A(n26), .ZN(N18) );
  INV_X1 U31 ( .A(n27), .ZN(N19) );
  INV_X1 U32 ( .A(n29), .ZN(N20) );
  INV_X1 U33 ( .A(n30), .ZN(N21) );
  INV_X1 U34 ( .A(n31), .ZN(N22) );
  INV_X1 U35 ( .A(n32), .ZN(N23) );
  INV_X1 U36 ( .A(n33), .ZN(N24) );
  INV_X1 U37 ( .A(n35), .ZN(N25) );
  INV_X1 U38 ( .A(n50), .ZN(N26) );
  INV_X1 U39 ( .A(n51), .ZN(N27) );
  INV_X1 U40 ( .A(n52), .ZN(N28) );
  INV_X1 U41 ( .A(n53), .ZN(N29) );
  INV_X1 U42 ( .A(n55), .ZN(N30) );
  INV_X1 U43 ( .A(n56), .ZN(N31) );
  INV_X1 U44 ( .A(n18), .ZN(N10) );
  INV_X1 U45 ( .A(n19), .ZN(N11) );
  INV_X1 U46 ( .A(n20), .ZN(N12) );
  AOI22_X1 U47 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U48 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U49 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U50 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U51 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U52 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U53 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U54 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U55 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U56 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U57 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U58 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U59 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U60 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U61 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U62 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U63 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U64 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U65 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U66 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_26 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n6), .Z(n17) );
  BUF_X1 U4 ( .A(n4), .Z(n9) );
  BUF_X1 U5 ( .A(n6), .Z(n15) );
  BUF_X1 U6 ( .A(n5), .Z(n14) );
  BUF_X1 U7 ( .A(n5), .Z(n12) );
  BUF_X1 U8 ( .A(n4), .Z(n11) );
  BUF_X1 U9 ( .A(n5), .Z(n13) );
  BUF_X1 U10 ( .A(n4), .Z(n10) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  AOI22_X1 U18 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U19 ( .A(n60), .ZN(N5) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U21 ( .A(n61), .ZN(N6) );
  AOI22_X1 U22 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U23 ( .A(n62), .ZN(N7) );
  AOI22_X1 U24 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U25 ( .A(n63), .ZN(N8) );
  AOI22_X1 U26 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n58), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U31 ( .A(n28), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U33 ( .A(n54), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U35 ( .A(n21), .ZN(N13) );
  AOI22_X1 U36 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U37 ( .A(n22), .ZN(N14) );
  AOI22_X1 U38 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U39 ( .A(n23), .ZN(N15) );
  AOI22_X1 U40 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U41 ( .A(n24), .ZN(N16) );
  AOI22_X1 U42 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U43 ( .A(n25), .ZN(N17) );
  AOI22_X1 U44 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U45 ( .A(n26), .ZN(N18) );
  AOI22_X1 U46 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U47 ( .A(n27), .ZN(N19) );
  AOI22_X1 U48 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U49 ( .A(n29), .ZN(N20) );
  AOI22_X1 U50 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U51 ( .A(n30), .ZN(N21) );
  AOI22_X1 U52 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U53 ( .A(n31), .ZN(N22) );
  AOI22_X1 U54 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U55 ( .A(n32), .ZN(N23) );
  AOI22_X1 U56 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U57 ( .A(n33), .ZN(N24) );
  AOI22_X1 U58 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U59 ( .A(n35), .ZN(N25) );
  AOI22_X1 U60 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U61 ( .A(n50), .ZN(N26) );
  AOI22_X1 U62 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U63 ( .A(n51), .ZN(N27) );
  AOI22_X1 U64 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U65 ( .A(n52), .ZN(N28) );
  AOI22_X1 U66 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U67 ( .A(n53), .ZN(N29) );
  AOI22_X1 U68 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U69 ( .A(n55), .ZN(N30) );
  AOI22_X1 U70 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U71 ( .A(n56), .ZN(N31) );
  AOI22_X1 U72 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U73 ( .A(n18), .ZN(N10) );
  AOI22_X1 U74 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U75 ( .A(n19), .ZN(N11) );
  AOI22_X1 U76 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U77 ( .A(n20), .ZN(N12) );
  AOI22_X1 U78 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_25 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n6), .Z(n17) );
  BUF_X1 U4 ( .A(n4), .Z(n9) );
  BUF_X1 U5 ( .A(n6), .Z(n15) );
  BUF_X1 U6 ( .A(n5), .Z(n14) );
  BUF_X1 U7 ( .A(n5), .Z(n12) );
  BUF_X1 U8 ( .A(n4), .Z(n11) );
  BUF_X1 U9 ( .A(n5), .Z(n13) );
  BUF_X1 U10 ( .A(n4), .Z(n10) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n64), .ZN(N9) );
  INV_X1 U16 ( .A(n59), .ZN(N4) );
  INV_X1 U17 ( .A(n60), .ZN(N5) );
  INV_X1 U18 ( .A(n61), .ZN(N6) );
  INV_X1 U19 ( .A(n62), .ZN(N7) );
  INV_X1 U20 ( .A(n63), .ZN(N8) );
  INV_X1 U21 ( .A(n57), .ZN(N32) );
  INV_X1 U22 ( .A(n58), .ZN(N33) );
  INV_X1 U23 ( .A(n28), .ZN(N2) );
  INV_X1 U24 ( .A(n54), .ZN(N3) );
  INV_X1 U25 ( .A(n21), .ZN(N13) );
  INV_X1 U26 ( .A(n22), .ZN(N14) );
  INV_X1 U27 ( .A(n23), .ZN(N15) );
  INV_X1 U28 ( .A(n24), .ZN(N16) );
  INV_X1 U29 ( .A(n25), .ZN(N17) );
  INV_X1 U30 ( .A(n26), .ZN(N18) );
  INV_X1 U31 ( .A(n27), .ZN(N19) );
  INV_X1 U32 ( .A(n29), .ZN(N20) );
  INV_X1 U33 ( .A(n30), .ZN(N21) );
  INV_X1 U34 ( .A(n31), .ZN(N22) );
  INV_X1 U35 ( .A(n32), .ZN(N23) );
  INV_X1 U36 ( .A(n33), .ZN(N24) );
  INV_X1 U37 ( .A(n35), .ZN(N25) );
  INV_X1 U38 ( .A(n50), .ZN(N26) );
  INV_X1 U39 ( .A(n51), .ZN(N27) );
  INV_X1 U40 ( .A(n52), .ZN(N28) );
  INV_X1 U41 ( .A(n53), .ZN(N29) );
  INV_X1 U42 ( .A(n55), .ZN(N30) );
  INV_X1 U43 ( .A(n56), .ZN(N31) );
  INV_X1 U44 ( .A(n18), .ZN(N10) );
  INV_X1 U45 ( .A(n19), .ZN(N11) );
  INV_X1 U46 ( .A(n20), .ZN(N12) );
  AOI22_X1 U47 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U48 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U49 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U50 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U51 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U52 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U53 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U54 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U55 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U56 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U57 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U58 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U59 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U60 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U61 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U62 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U63 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U64 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U65 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U66 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_24 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  INV_X1 U3 ( .A(n59), .ZN(N4) );
  INV_X1 U4 ( .A(n60), .ZN(N5) );
  INV_X1 U5 ( .A(n61), .ZN(N6) );
  INV_X1 U6 ( .A(n62), .ZN(N7) );
  INV_X1 U7 ( .A(n63), .ZN(N8) );
  INV_X1 U8 ( .A(n64), .ZN(N9) );
  INV_X1 U9 ( .A(n57), .ZN(N32) );
  INV_X1 U10 ( .A(n58), .ZN(N33) );
  INV_X1 U11 ( .A(n28), .ZN(N2) );
  INV_X1 U12 ( .A(n54), .ZN(N3) );
  INV_X1 U13 ( .A(n21), .ZN(N13) );
  INV_X1 U14 ( .A(n22), .ZN(N14) );
  INV_X1 U15 ( .A(n23), .ZN(N15) );
  INV_X1 U16 ( .A(n24), .ZN(N16) );
  INV_X1 U17 ( .A(n25), .ZN(N17) );
  INV_X1 U18 ( .A(n26), .ZN(N18) );
  INV_X1 U19 ( .A(n27), .ZN(N19) );
  INV_X1 U20 ( .A(n29), .ZN(N20) );
  INV_X1 U21 ( .A(n30), .ZN(N21) );
  INV_X1 U22 ( .A(n31), .ZN(N22) );
  INV_X1 U23 ( .A(n32), .ZN(N23) );
  INV_X1 U24 ( .A(n33), .ZN(N24) );
  INV_X1 U25 ( .A(n35), .ZN(N25) );
  INV_X1 U26 ( .A(n50), .ZN(N26) );
  INV_X1 U27 ( .A(n51), .ZN(N27) );
  INV_X1 U28 ( .A(n52), .ZN(N28) );
  INV_X1 U29 ( .A(n53), .ZN(N29) );
  INV_X1 U30 ( .A(n55), .ZN(N30) );
  INV_X1 U31 ( .A(n56), .ZN(N31) );
  INV_X1 U32 ( .A(n18), .ZN(N10) );
  INV_X1 U33 ( .A(n19), .ZN(N11) );
  INV_X1 U34 ( .A(n20), .ZN(N12) );
  BUF_X1 U35 ( .A(n4), .Z(n9) );
  BUF_X1 U36 ( .A(n6), .Z(n15) );
  BUF_X1 U37 ( .A(n5), .Z(n14) );
  BUF_X1 U38 ( .A(n5), .Z(n12) );
  BUF_X1 U39 ( .A(n4), .Z(n11) );
  BUF_X1 U40 ( .A(n5), .Z(n13) );
  BUF_X1 U41 ( .A(n4), .Z(n10) );
  BUF_X1 U42 ( .A(n6), .Z(n17) );
  BUF_X1 U43 ( .A(n6), .Z(n16) );
  AOI22_X1 U44 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U45 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U46 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U47 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U48 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U49 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U50 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U51 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U52 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U53 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U54 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U55 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U56 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U57 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U58 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U59 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U60 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U61 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U62 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U63 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U64 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U65 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U67 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U68 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U69 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U70 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U71 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U72 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  AOI22_X1 U73 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U74 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U75 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  BUF_X1 U76 ( .A(sel), .Z(n6) );
  BUF_X1 U77 ( .A(sel), .Z(n5) );
  BUF_X1 U78 ( .A(sel), .Z(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_23 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  INV_X1 U3 ( .A(n59), .ZN(N4) );
  INV_X1 U4 ( .A(n60), .ZN(N5) );
  INV_X1 U5 ( .A(n61), .ZN(N6) );
  INV_X1 U6 ( .A(n62), .ZN(N7) );
  INV_X1 U7 ( .A(n63), .ZN(N8) );
  INV_X1 U8 ( .A(n64), .ZN(N9) );
  INV_X1 U9 ( .A(n57), .ZN(N32) );
  INV_X1 U10 ( .A(n58), .ZN(N33) );
  INV_X1 U11 ( .A(n28), .ZN(N2) );
  INV_X1 U12 ( .A(n54), .ZN(N3) );
  INV_X1 U13 ( .A(n21), .ZN(N13) );
  INV_X1 U14 ( .A(n22), .ZN(N14) );
  INV_X1 U15 ( .A(n23), .ZN(N15) );
  INV_X1 U16 ( .A(n24), .ZN(N16) );
  INV_X1 U17 ( .A(n25), .ZN(N17) );
  INV_X1 U18 ( .A(n26), .ZN(N18) );
  INV_X1 U19 ( .A(n27), .ZN(N19) );
  INV_X1 U20 ( .A(n29), .ZN(N20) );
  INV_X1 U21 ( .A(n30), .ZN(N21) );
  INV_X1 U22 ( .A(n31), .ZN(N22) );
  INV_X1 U23 ( .A(n32), .ZN(N23) );
  INV_X1 U24 ( .A(n33), .ZN(N24) );
  INV_X1 U25 ( .A(n35), .ZN(N25) );
  INV_X1 U26 ( .A(n50), .ZN(N26) );
  INV_X1 U27 ( .A(n51), .ZN(N27) );
  INV_X1 U28 ( .A(n52), .ZN(N28) );
  INV_X1 U29 ( .A(n53), .ZN(N29) );
  INV_X1 U30 ( .A(n55), .ZN(N30) );
  INV_X1 U31 ( .A(n56), .ZN(N31) );
  INV_X1 U32 ( .A(n18), .ZN(N10) );
  INV_X1 U33 ( .A(n19), .ZN(N11) );
  INV_X1 U34 ( .A(n20), .ZN(N12) );
  BUF_X1 U35 ( .A(n4), .Z(n9) );
  BUF_X1 U36 ( .A(n6), .Z(n15) );
  BUF_X1 U37 ( .A(n5), .Z(n14) );
  BUF_X1 U38 ( .A(n5), .Z(n12) );
  BUF_X1 U39 ( .A(n4), .Z(n11) );
  BUF_X1 U40 ( .A(n5), .Z(n13) );
  BUF_X1 U41 ( .A(n4), .Z(n10) );
  BUF_X1 U42 ( .A(n6), .Z(n17) );
  BUF_X1 U43 ( .A(n6), .Z(n16) );
  AOI22_X1 U44 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U45 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U46 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U47 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U48 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U49 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U50 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U51 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U52 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U53 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U54 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U55 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U56 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U57 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U58 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U59 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U60 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U61 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U62 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U63 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U64 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U65 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U67 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U68 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U69 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U70 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U71 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U72 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  AOI22_X1 U73 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U74 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U75 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  BUF_X1 U76 ( .A(sel), .Z(n6) );
  BUF_X1 U77 ( .A(sel), .Z(n5) );
  BUF_X1 U78 ( .A(sel), .Z(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_22 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  INV_X1 U3 ( .A(n64), .ZN(N9) );
  INV_X1 U4 ( .A(n59), .ZN(N4) );
  INV_X1 U5 ( .A(n60), .ZN(N5) );
  INV_X1 U6 ( .A(n61), .ZN(N6) );
  INV_X1 U7 ( .A(n62), .ZN(N7) );
  INV_X1 U8 ( .A(n63), .ZN(N8) );
  INV_X1 U9 ( .A(n57), .ZN(N32) );
  INV_X1 U10 ( .A(n58), .ZN(N33) );
  INV_X1 U11 ( .A(n28), .ZN(N2) );
  INV_X1 U12 ( .A(n54), .ZN(N3) );
  INV_X1 U13 ( .A(n21), .ZN(N13) );
  INV_X1 U14 ( .A(n22), .ZN(N14) );
  INV_X1 U15 ( .A(n23), .ZN(N15) );
  INV_X1 U16 ( .A(n24), .ZN(N16) );
  INV_X1 U17 ( .A(n25), .ZN(N17) );
  INV_X1 U18 ( .A(n26), .ZN(N18) );
  INV_X1 U19 ( .A(n27), .ZN(N19) );
  INV_X1 U20 ( .A(n29), .ZN(N20) );
  INV_X1 U21 ( .A(n30), .ZN(N21) );
  INV_X1 U22 ( .A(n31), .ZN(N22) );
  INV_X1 U23 ( .A(n32), .ZN(N23) );
  INV_X1 U24 ( .A(n33), .ZN(N24) );
  INV_X1 U25 ( .A(n35), .ZN(N25) );
  INV_X1 U26 ( .A(n50), .ZN(N26) );
  INV_X1 U27 ( .A(n51), .ZN(N27) );
  INV_X1 U28 ( .A(n52), .ZN(N28) );
  INV_X1 U29 ( .A(n53), .ZN(N29) );
  INV_X1 U30 ( .A(n55), .ZN(N30) );
  INV_X1 U31 ( .A(n56), .ZN(N31) );
  INV_X1 U32 ( .A(n18), .ZN(N10) );
  INV_X1 U33 ( .A(n19), .ZN(N11) );
  INV_X1 U34 ( .A(n20), .ZN(N12) );
  BUF_X1 U35 ( .A(n4), .Z(n9) );
  BUF_X1 U36 ( .A(n6), .Z(n15) );
  BUF_X1 U37 ( .A(n5), .Z(n14) );
  BUF_X1 U38 ( .A(n5), .Z(n12) );
  BUF_X1 U39 ( .A(n4), .Z(n11) );
  BUF_X1 U40 ( .A(n5), .Z(n13) );
  BUF_X1 U41 ( .A(n4), .Z(n10) );
  BUF_X1 U42 ( .A(n6), .Z(n17) );
  BUF_X1 U43 ( .A(n6), .Z(n16) );
  AOI22_X1 U44 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U45 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U46 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U47 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U48 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U49 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U50 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U51 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U52 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U53 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U54 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U55 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U56 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U57 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U58 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U59 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U60 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U61 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U62 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U63 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U64 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U65 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U67 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U68 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U69 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U70 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U71 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U72 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  AOI22_X1 U73 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U74 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U75 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  BUF_X1 U76 ( .A(sel), .Z(n6) );
  BUF_X1 U77 ( .A(sel), .Z(n5) );
  BUF_X1 U78 ( .A(sel), .Z(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_21 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  INV_X1 U3 ( .A(n64), .ZN(N9) );
  INV_X1 U4 ( .A(n59), .ZN(N4) );
  INV_X1 U5 ( .A(n60), .ZN(N5) );
  INV_X1 U6 ( .A(n61), .ZN(N6) );
  INV_X1 U7 ( .A(n62), .ZN(N7) );
  INV_X1 U8 ( .A(n63), .ZN(N8) );
  INV_X1 U9 ( .A(n57), .ZN(N32) );
  INV_X1 U10 ( .A(n58), .ZN(N33) );
  INV_X1 U11 ( .A(n28), .ZN(N2) );
  INV_X1 U12 ( .A(n54), .ZN(N3) );
  INV_X1 U13 ( .A(n21), .ZN(N13) );
  INV_X1 U14 ( .A(n22), .ZN(N14) );
  INV_X1 U15 ( .A(n23), .ZN(N15) );
  INV_X1 U16 ( .A(n24), .ZN(N16) );
  INV_X1 U17 ( .A(n25), .ZN(N17) );
  INV_X1 U18 ( .A(n26), .ZN(N18) );
  INV_X1 U19 ( .A(n27), .ZN(N19) );
  INV_X1 U20 ( .A(n29), .ZN(N20) );
  INV_X1 U21 ( .A(n30), .ZN(N21) );
  INV_X1 U22 ( .A(n31), .ZN(N22) );
  INV_X1 U23 ( .A(n32), .ZN(N23) );
  INV_X1 U24 ( .A(n33), .ZN(N24) );
  INV_X1 U25 ( .A(n35), .ZN(N25) );
  INV_X1 U26 ( .A(n50), .ZN(N26) );
  INV_X1 U27 ( .A(n51), .ZN(N27) );
  INV_X1 U28 ( .A(n52), .ZN(N28) );
  INV_X1 U29 ( .A(n53), .ZN(N29) );
  INV_X1 U30 ( .A(n55), .ZN(N30) );
  INV_X1 U31 ( .A(n56), .ZN(N31) );
  INV_X1 U32 ( .A(n18), .ZN(N10) );
  INV_X1 U33 ( .A(n19), .ZN(N11) );
  INV_X1 U34 ( .A(n20), .ZN(N12) );
  BUF_X1 U35 ( .A(n4), .Z(n9) );
  BUF_X1 U36 ( .A(n6), .Z(n15) );
  BUF_X1 U37 ( .A(n5), .Z(n14) );
  BUF_X1 U38 ( .A(n5), .Z(n12) );
  BUF_X1 U39 ( .A(n4), .Z(n11) );
  BUF_X1 U40 ( .A(n5), .Z(n13) );
  BUF_X1 U41 ( .A(n4), .Z(n10) );
  BUF_X1 U42 ( .A(n6), .Z(n17) );
  BUF_X1 U43 ( .A(n6), .Z(n16) );
  AOI22_X1 U44 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U45 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U46 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U47 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U48 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U49 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U50 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U51 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U52 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U53 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U54 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U55 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U56 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U57 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U58 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U59 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U60 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U61 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U62 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U63 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U64 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U65 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U67 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U68 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U69 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U70 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U71 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U72 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  AOI22_X1 U73 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U74 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U75 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  BUF_X1 U76 ( .A(sel), .Z(n6) );
  BUF_X1 U77 ( .A(sel), .Z(n5) );
  BUF_X1 U78 ( .A(sel), .Z(n4) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_7 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  BUF_X1 U1 ( .A(sel), .Z(n5) );
  BUF_X1 U2 ( .A(n4), .Z(n11) );
  INV_X1 U3 ( .A(n35), .ZN(N28) );
  INV_X1 U4 ( .A(n49), .ZN(N30) );
  INV_X1 U5 ( .A(n47), .ZN(N29) );
  INV_X1 U6 ( .A(n50), .ZN(N31) );
  INV_X1 U7 ( .A(n33), .ZN(N27) );
  INV_X2 U8 ( .A(n5), .ZN(n8) );
  INV_X1 U9 ( .A(n10), .ZN(n7) );
  INV_X1 U10 ( .A(n32), .ZN(N26) );
  INV_X1 U11 ( .A(n31), .ZN(N25) );
  INV_X1 U12 ( .A(n29), .ZN(N23) );
  AOI22_X1 U13 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n29)
         );
  INV_X1 U14 ( .A(n30), .ZN(N24) );
  AOI22_X1 U15 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n30)
         );
  BUF_X1 U16 ( .A(n5), .Z(n13) );
  INV_X1 U17 ( .A(n23), .ZN(N18) );
  AOI22_X1 U18 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n23)
         );
  INV_X1 U19 ( .A(n28), .ZN(N22) );
  AOI22_X1 U20 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n28)
         );
  INV_X1 U21 ( .A(n22), .ZN(N17) );
  AOI22_X1 U22 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n22)
         );
  INV_X1 U23 ( .A(n26), .ZN(N20) );
  AOI22_X1 U24 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n26)
         );
  INV_X1 U25 ( .A(n24), .ZN(N19) );
  AOI22_X1 U26 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n24)
         );
  INV_X1 U27 ( .A(n27), .ZN(N21) );
  AOI22_X1 U28 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n27)
         );
  INV_X1 U29 ( .A(n20), .ZN(N15) );
  AOI22_X1 U30 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n14), .ZN(n20)
         );
  INV_X1 U31 ( .A(n19), .ZN(N14) );
  AOI22_X1 U32 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n14), .ZN(n19)
         );
  INV_X1 U33 ( .A(n17), .ZN(N12) );
  AOI22_X1 U34 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n14), .ZN(n17)
         );
  INV_X1 U35 ( .A(n21), .ZN(N16) );
  AOI22_X1 U36 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n14), .ZN(n21)
         );
  INV_X1 U37 ( .A(n18), .ZN(N13) );
  AOI22_X1 U38 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n14), .ZN(n18)
         );
  CLKBUF_X1 U39 ( .A(n5), .Z(n14) );
  CLKBUF_X1 U40 ( .A(n5), .Z(n12) );
  INV_X1 U41 ( .A(n16), .ZN(N11) );
  AOI22_X1 U42 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n14), .ZN(n16) );
  AOI22_X1 U43 ( .A1(port0[6]), .A2(n9), .B1(port1[6]), .B2(n10), .ZN(n57) );
  AOI22_X1 U44 ( .A1(port0[2]), .A2(n9), .B1(port1[2]), .B2(n14), .ZN(n53) );
  AOI22_X1 U45 ( .A1(port0[4]), .A2(n9), .B1(port1[4]), .B2(n10), .ZN(n55) );
  AOI22_X1 U46 ( .A1(port0[5]), .A2(n9), .B1(port1[5]), .B2(n10), .ZN(n56) );
  INV_X1 U47 ( .A(n57), .ZN(N8) );
  INV_X1 U48 ( .A(n53), .ZN(N4) );
  INV_X1 U49 ( .A(n55), .ZN(N6) );
  INV_X1 U50 ( .A(n56), .ZN(N7) );
  AOI22_X1 U51 ( .A1(port0[3]), .A2(n9), .B1(port1[3]), .B2(n10), .ZN(n54) );
  AOI22_X1 U52 ( .A1(port0[7]), .A2(n9), .B1(n14), .B2(port1[7]), .ZN(n58) );
  INV_X1 U53 ( .A(n54), .ZN(N5) );
  INV_X1 U54 ( .A(n58), .ZN(N9) );
  AOI22_X1 U55 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n25) );
  AOI22_X1 U56 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n48) );
  INV_X1 U57 ( .A(n25), .ZN(N2) );
  INV_X1 U58 ( .A(n48), .ZN(N3) );
  INV_X1 U59 ( .A(n15), .ZN(N10) );
  AOI22_X1 U60 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n14), .ZN(n15) );
  CLKBUF_X1 U61 ( .A(n4), .Z(n10) );
  CLKBUF_X1 U62 ( .A(sel), .Z(n6) );
  CLKBUF_X1 U63 ( .A(sel), .Z(n4) );
  AOI22_X1 U64 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n50)
         );
  AOI22_X1 U65 ( .A1(port0[30]), .A2(n9), .B1(port1[30]), .B2(n5), .ZN(n51) );
  AOI22_X1 U66 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n11), .ZN(n49)
         );
  AOI22_X1 U67 ( .A1(port0[31]), .A2(n9), .B1(port1[31]), .B2(n4), .ZN(n52) );
  INV_X1 U68 ( .A(n51), .ZN(N32) );
  AOI22_X1 U69 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n35)
         );
  AOI22_X1 U71 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n47)
         );
  INV_X1 U72 ( .A(n52), .ZN(N33) );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n33)
         );
  INV_X1 U75 ( .A(n6), .ZN(n9) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_6 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n44, n45, n46, n47, n48, n49, n50, n51, n52;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  BUF_X4 U1 ( .A(n5), .Z(n11) );
  BUF_X1 U2 ( .A(sel), .Z(n5) );
  BUF_X1 U3 ( .A(n4), .Z(n10) );
  INV_X1 U4 ( .A(n5), .ZN(n8) );
  INV_X1 U5 ( .A(n31), .ZN(N28) );
  INV_X1 U6 ( .A(n35), .ZN(N30) );
  INV_X1 U7 ( .A(n32), .ZN(N29) );
  INV_X1 U8 ( .A(n44), .ZN(N31) );
  INV_X1 U9 ( .A(n30), .ZN(N27) );
  INV_X1 U10 ( .A(n11), .ZN(n7) );
  INV_X1 U11 ( .A(n29), .ZN(N26) );
  AOI22_X1 U12 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n11), .ZN(n29)
         );
  AOI22_X1 U13 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n11), .ZN(n28)
         );
  INV_X1 U14 ( .A(n28), .ZN(N25) );
  INV_X1 U15 ( .A(n26), .ZN(N23) );
  INV_X1 U16 ( .A(n27), .ZN(N24) );
  INV_X1 U17 ( .A(n20), .ZN(N18) );
  INV_X1 U18 ( .A(n25), .ZN(N22) );
  INV_X1 U19 ( .A(n19), .ZN(N17) );
  INV_X1 U20 ( .A(n23), .ZN(N20) );
  INV_X1 U21 ( .A(n21), .ZN(N19) );
  INV_X1 U22 ( .A(n24), .ZN(N21) );
  AOI22_X1 U23 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n11), .ZN(n20)
         );
  AOI22_X1 U24 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n11), .ZN(n19)
         );
  AOI22_X1 U25 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n11), .ZN(n26)
         );
  AOI22_X1 U26 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n11), .ZN(n27)
         );
  AOI22_X1 U27 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n11), .ZN(n25)
         );
  AOI22_X1 U28 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n11), .ZN(n23)
         );
  AOI22_X1 U29 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n11), .ZN(n21)
         );
  AOI22_X1 U30 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n11), .ZN(n24)
         );
  AOI22_X1 U31 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n11), .ZN(n13) );
  AOI22_X1 U32 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n11), .ZN(n17)
         );
  AOI22_X1 U33 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n11), .ZN(n16)
         );
  AOI22_X1 U34 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n11), .ZN(n14)
         );
  AOI22_X1 U35 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n11), .ZN(n18)
         );
  INV_X1 U36 ( .A(n17), .ZN(N15) );
  INV_X1 U37 ( .A(n16), .ZN(N14) );
  INV_X1 U38 ( .A(n14), .ZN(N12) );
  INV_X1 U39 ( .A(n18), .ZN(N16) );
  AOI22_X1 U40 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n11), .ZN(n15)
         );
  INV_X1 U41 ( .A(n15), .ZN(N13) );
  INV_X1 U42 ( .A(n13), .ZN(N11) );
  INV_X1 U43 ( .A(n51), .ZN(N8) );
  INV_X1 U44 ( .A(n47), .ZN(N4) );
  INV_X1 U45 ( .A(n49), .ZN(N6) );
  INV_X1 U46 ( .A(n50), .ZN(N7) );
  INV_X1 U47 ( .A(n48), .ZN(N5) );
  INV_X1 U48 ( .A(n52), .ZN(N9) );
  AOI22_X1 U49 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n11), .ZN(n12) );
  INV_X1 U50 ( .A(n22), .ZN(N2) );
  AOI22_X1 U51 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n11), .ZN(n22) );
  INV_X1 U52 ( .A(n33), .ZN(N3) );
  AOI22_X1 U53 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n10), .ZN(n33) );
  INV_X1 U54 ( .A(n12), .ZN(N10) );
  CLKBUF_X1 U55 ( .A(sel), .Z(n6) );
  CLKBUF_X1 U56 ( .A(sel), .Z(n4) );
  AOI22_X1 U57 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n10), .ZN(n30)
         );
  INV_X1 U58 ( .A(n45), .ZN(N32) );
  AOI22_X1 U59 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n35)
         );
  AOI22_X1 U60 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n10), .ZN(n44)
         );
  AOI22_X1 U61 ( .A1(port0[2]), .A2(n9), .B1(port1[2]), .B2(n11), .ZN(n47) );
  AOI22_X1 U62 ( .A1(port0[3]), .A2(n9), .B1(port1[3]), .B2(n11), .ZN(n48) );
  AOI22_X1 U63 ( .A1(port0[4]), .A2(n9), .B1(port1[4]), .B2(n11), .ZN(n49) );
  AOI22_X1 U64 ( .A1(port0[5]), .A2(n9), .B1(port1[5]), .B2(n11), .ZN(n50) );
  AOI22_X1 U65 ( .A1(port0[6]), .A2(n9), .B1(port1[6]), .B2(n11), .ZN(n51) );
  AOI22_X1 U66 ( .A1(port0[7]), .A2(n9), .B1(n11), .B2(port1[7]), .ZN(n52) );
  AOI22_X1 U67 ( .A1(port0[30]), .A2(n9), .B1(port1[30]), .B2(n4), .ZN(n45) );
  AOI22_X1 U68 ( .A1(port0[31]), .A2(n9), .B1(port1[31]), .B2(n4), .ZN(n46) );
  INV_X1 U69 ( .A(n46), .ZN(N33) );
  AOI22_X1 U70 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n10), .ZN(n31)
         );
  AOI22_X1 U71 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n10), .ZN(n32)
         );
  INV_X1 U72 ( .A(n6), .ZN(n9) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_5 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  BUF_X2 U1 ( .A(n12), .Z(n8) );
  BUF_X1 U2 ( .A(n4), .Z(n12) );
  BUF_X1 U3 ( .A(sel), .Z(n13) );
  INV_X2 U4 ( .A(n13), .ZN(n6) );
  INV_X1 U5 ( .A(n33), .ZN(N28) );
  AOI22_X1 U6 ( .A1(port0[26]), .A2(n6), .B1(port1[26]), .B2(n12), .ZN(n33) );
  INV_X1 U7 ( .A(n47), .ZN(N30) );
  INV_X1 U8 ( .A(n32), .ZN(N27) );
  AOI22_X1 U9 ( .A1(port0[25]), .A2(n6), .B1(port1[25]), .B2(n8), .ZN(n32) );
  INV_X1 U10 ( .A(n48), .ZN(N31) );
  INV_X1 U11 ( .A(n35), .ZN(N29) );
  INV_X1 U12 ( .A(n13), .ZN(n5) );
  BUF_X1 U13 ( .A(n4), .Z(n11) );
  BUF_X1 U14 ( .A(sel), .Z(n9) );
  INV_X1 U15 ( .A(n22), .ZN(N18) );
  AOI22_X1 U16 ( .A1(port0[16]), .A2(n5), .B1(port1[16]), .B2(n12), .ZN(n22)
         );
  INV_X1 U17 ( .A(n27), .ZN(N22) );
  AOI22_X1 U18 ( .A1(port0[20]), .A2(n6), .B1(port1[20]), .B2(n11), .ZN(n27)
         );
  INV_X1 U19 ( .A(n21), .ZN(N17) );
  AOI22_X1 U20 ( .A1(port0[15]), .A2(n5), .B1(port1[15]), .B2(n12), .ZN(n21)
         );
  INV_X1 U21 ( .A(n25), .ZN(N20) );
  AOI22_X1 U22 ( .A1(port0[18]), .A2(n5), .B1(port1[18]), .B2(n11), .ZN(n25)
         );
  INV_X1 U23 ( .A(n23), .ZN(N19) );
  AOI22_X1 U24 ( .A1(port0[17]), .A2(n5), .B1(port1[17]), .B2(n12), .ZN(n23)
         );
  INV_X1 U25 ( .A(n26), .ZN(N21) );
  AOI22_X1 U26 ( .A1(port0[19]), .A2(n6), .B1(port1[19]), .B2(n11), .ZN(n26)
         );
  INV_X1 U27 ( .A(n16), .ZN(N12) );
  AOI22_X1 U28 ( .A1(port0[10]), .A2(n5), .B1(port1[10]), .B2(n8), .ZN(n16) );
  INV_X1 U29 ( .A(n20), .ZN(N16) );
  AOI22_X1 U30 ( .A1(port0[14]), .A2(n5), .B1(port1[14]), .B2(n8), .ZN(n20) );
  AOI22_X1 U31 ( .A1(port0[11]), .A2(n5), .B1(port1[11]), .B2(n8), .ZN(n17) );
  INV_X1 U32 ( .A(n17), .ZN(N13) );
  CLKBUF_X1 U33 ( .A(n4), .Z(n10) );
  INV_X1 U34 ( .A(n19), .ZN(N15) );
  AOI22_X1 U35 ( .A1(port0[13]), .A2(n5), .B1(port1[13]), .B2(n8), .ZN(n19) );
  INV_X1 U36 ( .A(n30), .ZN(N25) );
  AOI22_X1 U37 ( .A1(port0[23]), .A2(n6), .B1(port1[23]), .B2(n10), .ZN(n30)
         );
  INV_X1 U38 ( .A(n28), .ZN(N23) );
  AOI22_X1 U39 ( .A1(port0[21]), .A2(n6), .B1(port1[21]), .B2(n10), .ZN(n28)
         );
  INV_X1 U40 ( .A(n29), .ZN(N24) );
  AOI22_X1 U41 ( .A1(port0[22]), .A2(n6), .B1(port1[22]), .B2(n10), .ZN(n29)
         );
  INV_X1 U42 ( .A(n31), .ZN(N26) );
  AOI22_X1 U43 ( .A1(port0[24]), .A2(n6), .B1(port1[24]), .B2(n10), .ZN(n31)
         );
  INV_X1 U44 ( .A(n18), .ZN(N14) );
  AOI22_X1 U45 ( .A1(port0[12]), .A2(n5), .B1(port1[12]), .B2(n8), .ZN(n18) );
  INV_X1 U46 ( .A(n15), .ZN(N11) );
  AOI22_X1 U47 ( .A1(port0[9]), .A2(n5), .B1(port1[9]), .B2(n8), .ZN(n15) );
  AOI22_X1 U48 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n9), .ZN(n51) );
  AOI22_X1 U49 ( .A1(port0[4]), .A2(n7), .B1(port1[4]), .B2(n8), .ZN(n53) );
  AOI22_X1 U50 ( .A1(port0[5]), .A2(n7), .B1(port1[5]), .B2(n8), .ZN(n54) );
  INV_X1 U51 ( .A(n51), .ZN(N4) );
  INV_X1 U52 ( .A(n53), .ZN(N6) );
  INV_X1 U53 ( .A(n54), .ZN(N7) );
  AOI22_X1 U54 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n8), .ZN(n52) );
  INV_X1 U55 ( .A(n52), .ZN(N5) );
  AOI22_X1 U56 ( .A1(port0[1]), .A2(n6), .B1(port1[1]), .B2(n8), .ZN(n46) );
  INV_X1 U57 ( .A(n46), .ZN(N3) );
  INV_X1 U58 ( .A(n56), .ZN(N9) );
  AOI22_X1 U59 ( .A1(port0[7]), .A2(n7), .B1(n8), .B2(port1[7]), .ZN(n56) );
  INV_X1 U60 ( .A(n14), .ZN(N10) );
  AOI22_X1 U61 ( .A1(port0[8]), .A2(n5), .B1(port1[8]), .B2(n8), .ZN(n14) );
  INV_X1 U62 ( .A(n55), .ZN(N8) );
  AOI22_X1 U63 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n8), .ZN(n55) );
  INV_X1 U64 ( .A(n24), .ZN(N2) );
  AOI22_X1 U65 ( .A1(port0[0]), .A2(n5), .B1(port1[0]), .B2(n12), .ZN(n24) );
  CLKBUF_X1 U66 ( .A(sel), .Z(n4) );
  INV_X1 U67 ( .A(n49), .ZN(N32) );
  AOI22_X1 U68 ( .A1(port0[27]), .A2(n6), .B1(port1[27]), .B2(n10), .ZN(n35)
         );
  AOI22_X1 U69 ( .A1(port0[30]), .A2(n7), .B1(port1[30]), .B2(n9), .ZN(n49) );
  INV_X1 U70 ( .A(n50), .ZN(N33) );
  AOI22_X1 U71 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n9), .ZN(n50) );
  AOI22_X1 U72 ( .A1(port0[28]), .A2(n6), .B1(port1[28]), .B2(n9), .ZN(n47) );
  AOI22_X1 U73 ( .A1(port0[29]), .A2(n6), .B1(port1[29]), .B2(n11), .ZN(n48)
         );
  INV_X1 U74 ( .A(n13), .ZN(n7) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_4 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  BUF_X1 U1 ( .A(n10), .Z(n9) );
  BUF_X2 U2 ( .A(sel), .Z(n4) );
  INV_X1 U3 ( .A(n5), .ZN(n8) );
  INV_X2 U4 ( .A(n4), .ZN(n7) );
  INV_X1 U5 ( .A(n32), .ZN(N28) );
  INV_X1 U6 ( .A(n45), .ZN(N30) );
  INV_X1 U7 ( .A(n31), .ZN(N27) );
  AOI22_X1 U8 ( .A1(port0[28]), .A2(n7), .B1(port1[28]), .B2(n9), .ZN(n45) );
  AOI22_X1 U9 ( .A1(port0[27]), .A2(n7), .B1(port1[27]), .B2(n9), .ZN(n33) );
  INV_X1 U10 ( .A(n46), .ZN(N31) );
  INV_X1 U11 ( .A(n33), .ZN(N29) );
  INV_X1 U12 ( .A(n12), .ZN(n6) );
  AOI22_X1 U13 ( .A1(port0[26]), .A2(n7), .B1(port1[26]), .B2(n9), .ZN(n32) );
  AOI22_X1 U14 ( .A1(port0[25]), .A2(n7), .B1(port1[25]), .B2(n9), .ZN(n31) );
  BUF_X1 U15 ( .A(n4), .Z(n11) );
  INV_X1 U16 ( .A(n21), .ZN(N18) );
  INV_X1 U17 ( .A(n26), .ZN(N22) );
  INV_X1 U18 ( .A(n20), .ZN(N17) );
  INV_X1 U19 ( .A(n24), .ZN(N20) );
  INV_X1 U20 ( .A(n22), .ZN(N19) );
  INV_X1 U21 ( .A(n25), .ZN(N21) );
  AOI22_X1 U22 ( .A1(port0[16]), .A2(n6), .B1(port1[16]), .B2(n12), .ZN(n21)
         );
  AOI22_X1 U23 ( .A1(port0[23]), .A2(n7), .B1(port1[23]), .B2(n10), .ZN(n29)
         );
  AOI22_X1 U24 ( .A1(port0[15]), .A2(n6), .B1(port1[15]), .B2(n12), .ZN(n20)
         );
  AOI22_X1 U25 ( .A1(port0[21]), .A2(n7), .B1(port1[21]), .B2(n10), .ZN(n27)
         );
  AOI22_X1 U26 ( .A1(port0[22]), .A2(n7), .B1(port1[22]), .B2(n10), .ZN(n28)
         );
  AOI22_X1 U27 ( .A1(port0[20]), .A2(n7), .B1(port1[20]), .B2(n11), .ZN(n26)
         );
  AOI22_X1 U28 ( .A1(port0[24]), .A2(n7), .B1(port1[24]), .B2(n10), .ZN(n30)
         );
  AOI22_X1 U29 ( .A1(port0[17]), .A2(n6), .B1(port1[17]), .B2(n12), .ZN(n22)
         );
  AOI22_X1 U30 ( .A1(port0[18]), .A2(n6), .B1(port1[18]), .B2(n11), .ZN(n24)
         );
  AOI22_X1 U31 ( .A1(port0[19]), .A2(n7), .B1(port1[19]), .B2(n11), .ZN(n25)
         );
  AOI22_X1 U32 ( .A1(port0[9]), .A2(n6), .B1(port1[9]), .B2(n12), .ZN(n14) );
  AOI22_X1 U33 ( .A1(port0[13]), .A2(n6), .B1(port1[13]), .B2(n12), .ZN(n18)
         );
  AOI22_X1 U34 ( .A1(port0[12]), .A2(n6), .B1(port1[12]), .B2(n12), .ZN(n17)
         );
  AOI22_X1 U35 ( .A1(port0[10]), .A2(n6), .B1(port1[10]), .B2(n12), .ZN(n15)
         );
  AOI22_X1 U36 ( .A1(port0[14]), .A2(n6), .B1(port1[14]), .B2(n12), .ZN(n19)
         );
  INV_X1 U37 ( .A(n15), .ZN(N12) );
  INV_X1 U38 ( .A(n19), .ZN(N16) );
  INV_X1 U39 ( .A(n16), .ZN(N13) );
  AOI22_X1 U40 ( .A1(port0[11]), .A2(n6), .B1(port1[11]), .B2(n12), .ZN(n16)
         );
  CLKBUF_X1 U41 ( .A(n4), .Z(n12) );
  CLKBUF_X1 U42 ( .A(n4), .Z(n10) );
  INV_X1 U43 ( .A(n18), .ZN(N15) );
  INV_X1 U44 ( .A(n29), .ZN(N25) );
  INV_X1 U45 ( .A(n27), .ZN(N23) );
  INV_X1 U46 ( .A(n28), .ZN(N24) );
  INV_X1 U47 ( .A(n30), .ZN(N26) );
  INV_X1 U48 ( .A(n17), .ZN(N14) );
  INV_X1 U49 ( .A(n14), .ZN(N11) );
  INV_X1 U50 ( .A(n49), .ZN(N4) );
  AOI22_X1 U51 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n12), .ZN(n49) );
  INV_X1 U52 ( .A(n51), .ZN(N6) );
  AOI22_X1 U53 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n12), .ZN(n51) );
  INV_X1 U54 ( .A(n52), .ZN(N7) );
  AOI22_X1 U55 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n12), .ZN(n52) );
  INV_X1 U56 ( .A(n50), .ZN(N5) );
  AOI22_X1 U57 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n12), .ZN(n50) );
  AOI22_X1 U58 ( .A1(port0[7]), .A2(n8), .B1(n12), .B2(port1[7]), .ZN(n54) );
  AOI22_X1 U59 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n12), .ZN(n53) );
  AOI22_X1 U60 ( .A1(port0[8]), .A2(n6), .B1(port1[8]), .B2(n12), .ZN(n13) );
  INV_X1 U61 ( .A(n35), .ZN(N3) );
  AOI22_X1 U62 ( .A1(port0[1]), .A2(n7), .B1(port1[1]), .B2(n9), .ZN(n35) );
  INV_X1 U63 ( .A(n54), .ZN(N9) );
  INV_X1 U64 ( .A(n13), .ZN(N10) );
  INV_X1 U65 ( .A(n53), .ZN(N8) );
  INV_X1 U66 ( .A(n23), .ZN(N2) );
  CLKBUF_X1 U67 ( .A(sel), .Z(n5) );
  AOI22_X1 U68 ( .A1(port0[0]), .A2(n6), .B1(port1[0]), .B2(n12), .ZN(n23) );
  AOI22_X1 U69 ( .A1(port0[29]), .A2(n7), .B1(port1[29]), .B2(n11), .ZN(n46)
         );
  INV_X1 U70 ( .A(n47), .ZN(N32) );
  INV_X1 U71 ( .A(n48), .ZN(N33) );
  AOI22_X1 U72 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n4), .ZN(n47) );
  AOI22_X1 U73 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n4), .ZN(n48) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_137 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X2 U1 ( .A(n15), .ZN(n5) );
  BUF_X2 U2 ( .A(n3), .Z(n15) );
  INV_X2 U3 ( .A(n15), .ZN(n4) );
  CLKBUF_X1 U4 ( .A(n3), .Z(n14) );
  BUF_X1 U5 ( .A(n1), .Z(n8) );
  BUF_X1 U6 ( .A(n2), .Z(n10) );
  CLKBUF_X1 U7 ( .A(n1), .Z(n7) );
  BUF_X1 U8 ( .A(n2), .Z(n12) );
  CLKBUF_X1 U9 ( .A(n1), .Z(n9) );
  CLKBUF_X1 U10 ( .A(n2), .Z(n11) );
  BUF_X1 U11 ( .A(n3), .Z(n13) );
  BUF_X1 U12 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U13 ( .A(sel), .Z(n1) );
  CLKBUF_X1 U14 ( .A(sel), .Z(n2) );
  INV_X1 U15 ( .A(n53), .ZN(N32) );
  AOI22_X1 U16 ( .A1(port0[30]), .A2(n6), .B1(port1[30]), .B2(n8), .ZN(n53) );
  INV_X1 U17 ( .A(n58), .ZN(N7) );
  AOI22_X1 U18 ( .A1(port0[5]), .A2(n6), .B1(port1[5]), .B2(n7), .ZN(n58) );
  INV_X1 U19 ( .A(n55), .ZN(N4) );
  AOI22_X1 U20 ( .A1(port0[2]), .A2(n6), .B1(port1[2]), .B2(n8), .ZN(n55) );
  INV_X1 U21 ( .A(n31), .ZN(N24) );
  AOI22_X1 U22 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n10), .ZN(n31)
         );
  INV_X1 U23 ( .A(n32), .ZN(N25) );
  AOI22_X1 U24 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n10), .ZN(n32)
         );
  INV_X1 U25 ( .A(n51), .ZN(N30) );
  AOI22_X1 U26 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n8), .ZN(n51) );
  INV_X1 U27 ( .A(n29), .ZN(N22) );
  AOI22_X1 U28 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n11), .ZN(n29)
         );
  INV_X1 U29 ( .A(n28), .ZN(N21) );
  AOI22_X1 U30 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n11), .ZN(n28)
         );
  INV_X1 U31 ( .A(n27), .ZN(N20) );
  AOI22_X1 U32 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n11), .ZN(n27)
         );
  INV_X1 U33 ( .A(n57), .ZN(N6) );
  AOI22_X1 U34 ( .A1(port0[4]), .A2(n6), .B1(port1[4]), .B2(n7), .ZN(n57) );
  INV_X1 U35 ( .A(n59), .ZN(N8) );
  AOI22_X1 U36 ( .A1(port0[6]), .A2(n6), .B1(port1[6]), .B2(n7), .ZN(n59) );
  INV_X1 U37 ( .A(n60), .ZN(N9) );
  AOI22_X1 U38 ( .A1(port0[7]), .A2(n6), .B1(n14), .B2(port1[7]), .ZN(n60) );
  INV_X1 U39 ( .A(n21), .ZN(N15) );
  AOI22_X1 U40 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n13), .ZN(n21)
         );
  INV_X1 U41 ( .A(n16), .ZN(N10) );
  AOI22_X1 U42 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n14), .ZN(n16) );
  INV_X1 U43 ( .A(n19), .ZN(N13) );
  AOI22_X1 U44 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n13), .ZN(n19)
         );
  INV_X1 U45 ( .A(n24), .ZN(N18) );
  AOI22_X1 U46 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n12), .ZN(n24)
         );
  INV_X1 U47 ( .A(n25), .ZN(N19) );
  AOI22_X1 U48 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n12), .ZN(n25)
         );
  INV_X1 U49 ( .A(n26), .ZN(N2) );
  AOI22_X1 U50 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n12), .ZN(n26) );
  INV_X1 U51 ( .A(n56), .ZN(N5) );
  AOI22_X1 U52 ( .A1(port0[3]), .A2(n6), .B1(port1[3]), .B2(n7), .ZN(n56) );
  INV_X1 U53 ( .A(n54), .ZN(N33) );
  AOI22_X1 U54 ( .A1(port0[31]), .A2(n6), .B1(port1[31]), .B2(n8), .ZN(n54) );
  INV_X1 U55 ( .A(n48), .ZN(N28) );
  AOI22_X1 U56 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n9), .ZN(n48) );
  INV_X1 U57 ( .A(n50), .ZN(N3) );
  AOI22_X1 U58 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n9), .ZN(n50) );
  INV_X1 U59 ( .A(n30), .ZN(N23) );
  AOI22_X1 U60 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n10), .ZN(n30)
         );
  INV_X1 U61 ( .A(n52), .ZN(N31) );
  AOI22_X1 U62 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n11), .ZN(n52)
         );
  INV_X1 U63 ( .A(n22), .ZN(N16) );
  AOI22_X1 U64 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n13), .ZN(n22)
         );
  INV_X1 U65 ( .A(n23), .ZN(N17) );
  AOI22_X1 U66 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n12), .ZN(n23)
         );
  INV_X1 U67 ( .A(n20), .ZN(N14) );
  AOI22_X1 U68 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n13), .ZN(n20)
         );
  INV_X1 U69 ( .A(n18), .ZN(N12) );
  AOI22_X1 U70 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n14), .ZN(n18)
         );
  INV_X1 U71 ( .A(n49), .ZN(N29) );
  AOI22_X1 U72 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n9), .ZN(n49) );
  INV_X1 U73 ( .A(n17), .ZN(N11) );
  AOI22_X1 U74 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n14), .ZN(n17) );
  INV_X1 U75 ( .A(n33), .ZN(N26) );
  AOI22_X1 U76 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n10), .ZN(n33)
         );
  INV_X1 U77 ( .A(n35), .ZN(N27) );
  AOI22_X1 U78 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n9), .ZN(n35) );
  INV_X1 U79 ( .A(n15), .ZN(n6) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_136 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  BUF_X1 U1 ( .A(n3), .Z(n9) );
  CLKBUF_X1 U2 ( .A(n3), .Z(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n15) );
  BUF_X2 U4 ( .A(n14), .Z(n10) );
  CLKBUF_X1 U5 ( .A(n3), .Z(n11) );
  BUF_X1 U6 ( .A(n3), .Z(n12) );
  BUF_X2 U7 ( .A(n3), .Z(n14) );
  BUF_X2 U8 ( .A(sel), .Z(n3) );
  INV_X1 U9 ( .A(n15), .ZN(n1) );
  INV_X1 U10 ( .A(n15), .ZN(n6) );
  CLKBUF_X1 U11 ( .A(n3), .Z(n13) );
  INV_X1 U12 ( .A(n4), .ZN(n5) );
  INV_X1 U13 ( .A(n53), .ZN(N32) );
  INV_X1 U14 ( .A(n58), .ZN(N7) );
  INV_X1 U15 ( .A(n31), .ZN(N24) );
  INV_X1 U16 ( .A(n32), .ZN(N25) );
  INV_X1 U17 ( .A(n28), .ZN(N21) );
  INV_X1 U18 ( .A(n16), .ZN(N10) );
  INV_X1 U19 ( .A(n20), .ZN(N14) );
  INV_X1 U20 ( .A(n19), .ZN(N13) );
  INV_X1 U21 ( .A(n49), .ZN(N29) );
  INV_X1 U22 ( .A(n33), .ZN(N26) );
  INV_X1 U23 ( .A(n50), .ZN(N3) );
  INV_X1 U24 ( .A(n27), .ZN(N20) );
  INV_X1 U25 ( .A(n25), .ZN(N19) );
  INV_X1 U26 ( .A(n35), .ZN(N27) );
  INV_X1 U27 ( .A(n60), .ZN(N9) );
  INV_X1 U28 ( .A(n59), .ZN(N8) );
  INV_X1 U29 ( .A(n55), .ZN(N4) );
  INV_X1 U30 ( .A(n56), .ZN(N5) );
  INV_X1 U31 ( .A(n48), .ZN(N28) );
  INV_X1 U32 ( .A(n30), .ZN(N23) );
  INV_X1 U33 ( .A(n52), .ZN(N31) );
  INV_X1 U34 ( .A(n22), .ZN(N16) );
  INV_X1 U35 ( .A(n51), .ZN(N30) );
  INV_X1 U36 ( .A(n29), .ZN(N22) );
  INV_X1 U37 ( .A(n23), .ZN(N17) );
  INV_X1 U38 ( .A(n21), .ZN(N15) );
  INV_X1 U39 ( .A(n18), .ZN(N12) );
  INV_X1 U40 ( .A(n17), .ZN(N11) );
  INV_X1 U41 ( .A(n24), .ZN(N18) );
  INV_X1 U42 ( .A(n26), .ZN(N2) );
  INV_X1 U43 ( .A(n57), .ZN(N6) );
  AOI22_X1 U44 ( .A1(port0[26]), .A2(n1), .B1(port1[26]), .B2(n9), .ZN(n48) );
  AOI22_X1 U45 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n10), .ZN(n31)
         );
  AOI22_X1 U46 ( .A1(port0[21]), .A2(n1), .B1(port1[21]), .B2(n10), .ZN(n30)
         );
  AOI22_X1 U47 ( .A1(port0[29]), .A2(n6), .B1(port1[29]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n1), .B1(port1[14]), .B2(n13), .ZN(n22)
         );
  AOI22_X1 U49 ( .A1(port0[23]), .A2(n6), .B1(port1[23]), .B2(n10), .ZN(n32)
         );
  AOI22_X1 U50 ( .A1(port0[28]), .A2(n2), .B1(port1[28]), .B2(n8), .ZN(n51) );
  AOI22_X1 U51 ( .A1(port0[20]), .A2(n1), .B1(port1[20]), .B2(n11), .ZN(n29)
         );
  AOI22_X1 U52 ( .A1(port0[15]), .A2(n6), .B1(port1[15]), .B2(n12), .ZN(n23)
         );
  AOI22_X1 U53 ( .A1(port0[13]), .A2(n1), .B1(port1[13]), .B2(n13), .ZN(n21)
         );
  AOI22_X1 U54 ( .A1(port0[19]), .A2(n1), .B1(port1[19]), .B2(n11), .ZN(n28)
         );
  AOI22_X1 U55 ( .A1(port0[8]), .A2(n6), .B1(port1[8]), .B2(n14), .ZN(n16) );
  AOI22_X1 U56 ( .A1(port0[12]), .A2(n5), .B1(port1[12]), .B2(n13), .ZN(n20)
         );
  AOI22_X1 U57 ( .A1(port0[10]), .A2(n1), .B1(port1[10]), .B2(n14), .ZN(n18)
         );
  AOI22_X1 U58 ( .A1(port0[11]), .A2(n1), .B1(port1[11]), .B2(n13), .ZN(n19)
         );
  AOI22_X1 U59 ( .A1(port0[27]), .A2(n6), .B1(port1[27]), .B2(n9), .ZN(n49) );
  AOI22_X1 U60 ( .A1(port0[9]), .A2(n2), .B1(port1[9]), .B2(n14), .ZN(n17) );
  AOI22_X1 U61 ( .A1(port0[24]), .A2(n1), .B1(port1[24]), .B2(n10), .ZN(n33)
         );
  AOI22_X1 U62 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n9), .ZN(n50) );
  AOI22_X1 U63 ( .A1(port0[18]), .A2(n1), .B1(port1[18]), .B2(n11), .ZN(n27)
         );
  AOI22_X1 U64 ( .A1(port0[16]), .A2(n1), .B1(port1[16]), .B2(n12), .ZN(n24)
         );
  AOI22_X1 U65 ( .A1(port0[17]), .A2(n1), .B1(port1[17]), .B2(n12), .ZN(n25)
         );
  AOI22_X1 U66 ( .A1(port0[25]), .A2(n6), .B1(port1[25]), .B2(n9), .ZN(n35) );
  AOI22_X1 U67 ( .A1(port0[0]), .A2(n5), .B1(port1[0]), .B2(n12), .ZN(n26) );
  INV_X1 U68 ( .A(n3), .ZN(n2) );
  CLKBUF_X1 U69 ( .A(n3), .Z(n7) );
  BUF_X1 U70 ( .A(sel), .Z(n4) );
  AOI22_X1 U71 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n8), .ZN(n53) );
  AOI22_X1 U72 ( .A1(port0[2]), .A2(n2), .B1(port1[2]), .B2(n8), .ZN(n55) );
  AOI22_X1 U73 ( .A1(port0[7]), .A2(n2), .B1(n14), .B2(port1[7]), .ZN(n60) );
  AOI22_X1 U74 ( .A1(port0[5]), .A2(n2), .B1(port1[5]), .B2(n7), .ZN(n58) );
  AOI22_X1 U75 ( .A1(port0[3]), .A2(n2), .B1(port1[3]), .B2(n7), .ZN(n56) );
  AOI22_X1 U76 ( .A1(port0[4]), .A2(n2), .B1(port1[4]), .B2(n7), .ZN(n57) );
  AOI22_X1 U77 ( .A1(port0[6]), .A2(n2), .B1(port1[6]), .B2(n7), .ZN(n59) );
  INV_X1 U78 ( .A(n54), .ZN(N33) );
  AOI22_X1 U79 ( .A1(n5), .A2(port0[31]), .B1(port1[31]), .B2(n8), .ZN(n54) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_135 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N32, N33, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n35, n43, n51, n52, n53, n54, n55, n56, n57,
         n58, n59, n60, n61, n62, n63, n64, n65;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[30] = N32;
  assign portY[31] = N33;

  CLKBUF_X1 U1 ( .A(n7), .Z(n19) );
  CLKBUF_X1 U2 ( .A(n5), .Z(n13) );
  BUF_X2 U3 ( .A(n5), .Z(n12) );
  CLKBUF_X1 U4 ( .A(n5), .Z(n11) );
  BUF_X2 U5 ( .A(sel), .Z(n7) );
  NAND2_X1 U6 ( .A1(port0[29]), .A2(n9), .ZN(n1) );
  NAND2_X1 U7 ( .A1(port1[29]), .A2(n15), .ZN(n2) );
  NAND2_X1 U8 ( .A1(n1), .A2(n2), .ZN(portY[29]) );
  CLKBUF_X1 U9 ( .A(sel), .Z(n5) );
  BUF_X1 U10 ( .A(n6), .Z(n15) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  INV_X2 U12 ( .A(n7), .ZN(n10) );
  INV_X1 U13 ( .A(n19), .ZN(n8) );
  INV_X1 U14 ( .A(n5), .ZN(n4) );
  INV_X1 U15 ( .A(n7), .ZN(n9) );
  CLKBUF_X1 U16 ( .A(n6), .Z(n17) );
  CLKBUF_X1 U17 ( .A(n5), .Z(n14) );
  INV_X1 U18 ( .A(n58), .ZN(N32) );
  INV_X1 U19 ( .A(n63), .ZN(N7) );
  INV_X1 U20 ( .A(n43), .ZN(N24) );
  INV_X1 U21 ( .A(n51), .ZN(N25) );
  INV_X1 U22 ( .A(n32), .ZN(N21) );
  INV_X1 U23 ( .A(n20), .ZN(N10) );
  INV_X1 U24 ( .A(n24), .ZN(N14) );
  INV_X1 U25 ( .A(n23), .ZN(N13) );
  INV_X1 U26 ( .A(n55), .ZN(N29) );
  INV_X1 U27 ( .A(n52), .ZN(N26) );
  INV_X1 U28 ( .A(n56), .ZN(N3) );
  INV_X1 U29 ( .A(n31), .ZN(N20) );
  INV_X1 U30 ( .A(n29), .ZN(N19) );
  INV_X1 U31 ( .A(n53), .ZN(N27) );
  INV_X1 U32 ( .A(n65), .ZN(N9) );
  INV_X1 U33 ( .A(n64), .ZN(N8) );
  INV_X1 U34 ( .A(n60), .ZN(N4) );
  INV_X1 U35 ( .A(n61), .ZN(N5) );
  INV_X1 U36 ( .A(n54), .ZN(N28) );
  INV_X1 U37 ( .A(n35), .ZN(N23) );
  INV_X1 U38 ( .A(n26), .ZN(N16) );
  INV_X1 U39 ( .A(n57), .ZN(N30) );
  INV_X1 U40 ( .A(n33), .ZN(N22) );
  INV_X1 U41 ( .A(n27), .ZN(N17) );
  INV_X1 U42 ( .A(n25), .ZN(N15) );
  INV_X1 U43 ( .A(n22), .ZN(N12) );
  INV_X1 U44 ( .A(n21), .ZN(N11) );
  INV_X1 U45 ( .A(n28), .ZN(N18) );
  INV_X1 U46 ( .A(n30), .ZN(N2) );
  INV_X1 U47 ( .A(n62), .ZN(N6) );
  AOI22_X1 U48 ( .A1(port0[26]), .A2(n10), .B1(port1[26]), .B2(n12), .ZN(n54)
         );
  AOI22_X1 U49 ( .A1(port0[22]), .A2(n10), .B1(port1[22]), .B2(n11), .ZN(n43)
         );
  AOI22_X1 U50 ( .A1(port0[21]), .A2(n10), .B1(port1[21]), .B2(n11), .ZN(n35)
         );
  AOI22_X1 U51 ( .A1(port0[23]), .A2(n10), .B1(port1[23]), .B2(n14), .ZN(n51)
         );
  AOI22_X1 U52 ( .A1(port0[28]), .A2(n9), .B1(port1[28]), .B2(n14), .ZN(n57)
         );
  AOI22_X1 U53 ( .A1(port0[20]), .A2(n10), .B1(port1[20]), .B2(n15), .ZN(n33)
         );
  AOI22_X1 U54 ( .A1(port0[19]), .A2(n10), .B1(port1[19]), .B2(n15), .ZN(n32)
         );
  AOI22_X1 U55 ( .A1(port0[27]), .A2(n10), .B1(port1[27]), .B2(n12), .ZN(n55)
         );
  AOI22_X1 U56 ( .A1(port0[24]), .A2(n10), .B1(port1[24]), .B2(n12), .ZN(n52)
         );
  AOI22_X1 U57 ( .A1(port0[1]), .A2(n9), .B1(port1[1]), .B2(n13), .ZN(n56) );
  AOI22_X1 U58 ( .A1(port0[25]), .A2(n10), .B1(port1[25]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U59 ( .A1(port0[8]), .A2(n8), .B1(port1[8]), .B2(n18), .ZN(n20) );
  AOI22_X1 U60 ( .A1(port0[9]), .A2(n8), .B1(port1[9]), .B2(n18), .ZN(n21) );
  AOI22_X1 U61 ( .A1(port0[10]), .A2(n8), .B1(port1[10]), .B2(n18), .ZN(n22)
         );
  AOI22_X1 U62 ( .A1(port0[11]), .A2(n8), .B1(port1[11]), .B2(n17), .ZN(n23)
         );
  AOI22_X1 U63 ( .A1(port0[12]), .A2(n8), .B1(port1[12]), .B2(n17), .ZN(n24)
         );
  AOI22_X1 U64 ( .A1(port0[13]), .A2(n8), .B1(port1[13]), .B2(n17), .ZN(n25)
         );
  AOI22_X1 U65 ( .A1(port0[14]), .A2(n8), .B1(port1[14]), .B2(n17), .ZN(n26)
         );
  AOI22_X1 U66 ( .A1(port0[15]), .A2(n8), .B1(port1[15]), .B2(n16), .ZN(n27)
         );
  AOI22_X1 U67 ( .A1(port0[16]), .A2(n8), .B1(port1[16]), .B2(n16), .ZN(n28)
         );
  AOI22_X1 U68 ( .A1(port0[17]), .A2(n8), .B1(port1[17]), .B2(n16), .ZN(n29)
         );
  AOI22_X1 U69 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n16), .ZN(n30) );
  AOI22_X1 U70 ( .A1(port0[18]), .A2(n8), .B1(port1[18]), .B2(n15), .ZN(n31)
         );
  CLKBUF_X1 U71 ( .A(n6), .Z(n18) );
  CLKBUF_X1 U72 ( .A(sel), .Z(n6) );
  AOI22_X1 U73 ( .A1(port0[2]), .A2(n10), .B1(port1[2]), .B2(n14), .ZN(n60) );
  AOI22_X1 U74 ( .A1(port0[5]), .A2(n10), .B1(port1[5]), .B2(n12), .ZN(n63) );
  AOI22_X1 U75 ( .A1(port0[4]), .A2(n10), .B1(port1[4]), .B2(n14), .ZN(n62) );
  AOI22_X1 U76 ( .A1(port0[3]), .A2(n10), .B1(port1[3]), .B2(n12), .ZN(n61) );
  AOI22_X1 U77 ( .A1(port0[7]), .A2(n10), .B1(n18), .B2(port1[7]), .ZN(n65) );
  AOI22_X1 U78 ( .A1(port0[6]), .A2(n10), .B1(port1[6]), .B2(n11), .ZN(n64) );
  AOI22_X1 U79 ( .A1(port0[30]), .A2(n9), .B1(port1[30]), .B2(n13), .ZN(n58)
         );
  AOI22_X1 U80 ( .A1(port0[31]), .A2(n9), .B1(port1[31]), .B2(n11), .ZN(n59)
         );
  INV_X1 U81 ( .A(n59), .ZN(N33) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_134 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n41, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  MUX2_X1 U1 ( .A(port0[0]), .B(port1[0]), .S(sel), .Z(N2) );
  MUX2_X1 U2 ( .A(port0[31]), .B(port1[31]), .S(sel), .Z(N33) );
  BUF_X2 U3 ( .A(n5), .Z(n17) );
  BUF_X1 U4 ( .A(sel), .Z(n3) );
  BUF_X1 U5 ( .A(sel), .Z(n4) );
  INV_X1 U6 ( .A(n17), .ZN(n1) );
  INV_X1 U7 ( .A(n17), .ZN(n7) );
  INV_X1 U8 ( .A(n17), .ZN(n2) );
  INV_X1 U9 ( .A(n17), .ZN(n6) );
  BUF_X1 U10 ( .A(n4), .Z(n14) );
  CLKBUF_X1 U11 ( .A(n3), .Z(n11) );
  CLKBUF_X1 U12 ( .A(n5), .Z(n15) );
  CLKBUF_X1 U13 ( .A(n5), .Z(n16) );
  BUF_X1 U14 ( .A(n4), .Z(n12) );
  CLKBUF_X1 U15 ( .A(n4), .Z(n13) );
  BUF_X1 U16 ( .A(n3), .Z(n10) );
  CLKBUF_X1 U17 ( .A(n3), .Z(n9) );
  BUF_X1 U18 ( .A(sel), .Z(n5) );
  INV_X1 U19 ( .A(n57), .ZN(N7) );
  INV_X1 U20 ( .A(n32), .ZN(N24) );
  AOI22_X1 U21 ( .A1(port0[22]), .A2(n2), .B1(port1[22]), .B2(n12), .ZN(n32)
         );
  INV_X1 U22 ( .A(n33), .ZN(N25) );
  AOI22_X1 U23 ( .A1(port0[23]), .A2(n6), .B1(port1[23]), .B2(n12), .ZN(n33)
         );
  INV_X1 U24 ( .A(n29), .ZN(N21) );
  AOI22_X1 U25 ( .A1(port0[19]), .A2(n2), .B1(port1[19]), .B2(n13), .ZN(n29)
         );
  INV_X1 U26 ( .A(n18), .ZN(N10) );
  AOI22_X1 U27 ( .A1(port0[8]), .A2(n1), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U28 ( .A(n22), .ZN(N14) );
  AOI22_X1 U29 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U30 ( .A(n21), .ZN(N13) );
  AOI22_X1 U31 ( .A1(port0[11]), .A2(n2), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U32 ( .A(n49), .ZN(N29) );
  AOI22_X1 U33 ( .A1(port0[27]), .A2(n2), .B1(port1[27]), .B2(n11), .ZN(n49)
         );
  INV_X1 U34 ( .A(n35), .ZN(N26) );
  AOI22_X1 U35 ( .A1(port0[24]), .A2(n6), .B1(port1[24]), .B2(n12), .ZN(n35)
         );
  INV_X1 U36 ( .A(n50), .ZN(N3) );
  AOI22_X1 U37 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n50) );
  INV_X1 U38 ( .A(n28), .ZN(N20) );
  AOI22_X1 U39 ( .A1(port0[18]), .A2(n6), .B1(port1[18]), .B2(n13), .ZN(n28)
         );
  INV_X1 U40 ( .A(n27), .ZN(N19) );
  AOI22_X1 U41 ( .A1(port0[17]), .A2(n1), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U42 ( .A(n41), .ZN(N27) );
  AOI22_X1 U43 ( .A1(port0[25]), .A2(n7), .B1(port1[25]), .B2(n11), .ZN(n41)
         );
  INV_X1 U44 ( .A(n59), .ZN(N9) );
  INV_X1 U45 ( .A(n58), .ZN(N8) );
  INV_X1 U46 ( .A(n54), .ZN(N4) );
  INV_X1 U47 ( .A(n55), .ZN(N5) );
  INV_X1 U48 ( .A(n48), .ZN(N28) );
  AOI22_X1 U49 ( .A1(port0[26]), .A2(n6), .B1(port1[26]), .B2(n11), .ZN(n48)
         );
  INV_X1 U50 ( .A(n31), .ZN(N23) );
  AOI22_X1 U51 ( .A1(port0[21]), .A2(n1), .B1(port1[21]), .B2(n12), .ZN(n31)
         );
  INV_X1 U52 ( .A(n52), .ZN(N31) );
  AOI22_X1 U53 ( .A1(port0[29]), .A2(n1), .B1(port1[29]), .B2(n13), .ZN(n52)
         );
  INV_X1 U54 ( .A(n24), .ZN(N16) );
  AOI22_X1 U55 ( .A1(port0[14]), .A2(n6), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U56 ( .A(n51), .ZN(N30) );
  AOI22_X1 U57 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n51)
         );
  INV_X1 U58 ( .A(n30), .ZN(N22) );
  AOI22_X1 U59 ( .A1(port0[20]), .A2(n7), .B1(port1[20]), .B2(n13), .ZN(n30)
         );
  INV_X1 U60 ( .A(n25), .ZN(N17) );
  AOI22_X1 U61 ( .A1(port0[15]), .A2(n2), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U62 ( .A(n23), .ZN(N15) );
  AOI22_X1 U63 ( .A1(port0[13]), .A2(n2), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U64 ( .A(n20), .ZN(N12) );
  AOI22_X1 U65 ( .A1(port0[10]), .A2(n1), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U66 ( .A(n19), .ZN(N11) );
  AOI22_X1 U67 ( .A1(port0[9]), .A2(n6), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U68 ( .A(n26), .ZN(N18) );
  AOI22_X1 U69 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U70 ( .A(n56), .ZN(N6) );
  INV_X1 U71 ( .A(n17), .ZN(n8) );
  AOI22_X1 U72 ( .A1(port0[2]), .A2(n1), .B1(port1[2]), .B2(n10), .ZN(n54) );
  AOI22_X1 U73 ( .A1(port0[5]), .A2(n6), .B1(port1[5]), .B2(n9), .ZN(n57) );
  AOI22_X1 U74 ( .A1(port0[7]), .A2(n6), .B1(n16), .B2(port1[7]), .ZN(n59) );
  AOI22_X1 U75 ( .A1(port0[4]), .A2(n6), .B1(port1[4]), .B2(n9), .ZN(n56) );
  AOI22_X1 U76 ( .A1(port0[3]), .A2(n6), .B1(port1[3]), .B2(n9), .ZN(n55) );
  AOI22_X1 U77 ( .A1(port0[6]), .A2(n7), .B1(port1[6]), .B2(n9), .ZN(n58) );
  AOI22_X1 U78 ( .A1(n7), .A2(port0[30]), .B1(port1[30]), .B2(n10), .ZN(n53)
         );
  INV_X1 U79 ( .A(n53), .ZN(N32) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_133 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  CLKBUF_X3 U1 ( .A(n11), .Z(n5) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n8) );
  BUF_X1 U3 ( .A(sel), .Z(n9) );
  INV_X1 U4 ( .A(n7), .ZN(n1) );
  BUF_X1 U5 ( .A(sel), .Z(n7) );
  BUF_X2 U6 ( .A(n9), .Z(n15) );
  BUF_X1 U7 ( .A(n10), .Z(n6) );
  INV_X1 U8 ( .A(n12), .ZN(n2) );
  BUF_X2 U9 ( .A(n7), .Z(n12) );
  BUF_X2 U10 ( .A(n9), .Z(n13) );
  INV_X1 U11 ( .A(n15), .ZN(n3) );
  BUF_X1 U12 ( .A(n10), .Z(n4) );
  INV_X1 U13 ( .A(n9), .ZN(n10) );
  CLKBUF_X1 U14 ( .A(n8), .Z(n14) );
  INV_X1 U15 ( .A(n7), .ZN(n11) );
  INV_X1 U16 ( .A(n50), .ZN(N3) );
  INV_X1 U17 ( .A(n33), .ZN(N26) );
  INV_X1 U18 ( .A(n57), .ZN(N6) );
  INV_X1 U19 ( .A(n55), .ZN(N4) );
  INV_X1 U20 ( .A(n53), .ZN(N32) );
  INV_X1 U21 ( .A(n26), .ZN(N2) );
  INV_X1 U22 ( .A(n60), .ZN(N9) );
  INV_X1 U23 ( .A(n58), .ZN(N7) );
  INV_X1 U24 ( .A(n31), .ZN(N24) );
  INV_X1 U25 ( .A(n30), .ZN(N23) );
  INV_X1 U26 ( .A(n32), .ZN(N25) );
  INV_X1 U27 ( .A(n23), .ZN(N17) );
  INV_X1 U28 ( .A(n28), .ZN(N21) );
  INV_X1 U29 ( .A(n16), .ZN(N10) );
  INV_X1 U30 ( .A(n20), .ZN(N14) );
  INV_X1 U31 ( .A(n19), .ZN(N13) );
  INV_X1 U32 ( .A(n49), .ZN(N29) );
  INV_X1 U33 ( .A(n35), .ZN(N27) );
  INV_X1 U34 ( .A(n48), .ZN(N28) );
  INV_X1 U35 ( .A(n52), .ZN(N31) );
  INV_X1 U36 ( .A(n22), .ZN(N16) );
  INV_X1 U37 ( .A(n59), .ZN(N8) );
  INV_X1 U38 ( .A(n29), .ZN(N22) );
  INV_X1 U39 ( .A(n51), .ZN(N30) );
  INV_X1 U40 ( .A(n21), .ZN(N15) );
  INV_X1 U41 ( .A(n18), .ZN(N12) );
  INV_X1 U42 ( .A(n17), .ZN(N11) );
  INV_X1 U43 ( .A(n27), .ZN(N20) );
  INV_X1 U44 ( .A(n24), .ZN(N18) );
  INV_X1 U45 ( .A(n25), .ZN(N19) );
  AOI22_X1 U46 ( .A1(port0[26]), .A2(n1), .B1(port1[26]), .B2(n15), .ZN(n48)
         );
  AOI22_X1 U47 ( .A1(port0[1]), .A2(n10), .B1(port1[1]), .B2(n8), .ZN(n50) );
  AOI22_X1 U48 ( .A1(port0[21]), .A2(n3), .B1(port1[21]), .B2(n12), .ZN(n30)
         );
  AOI22_X1 U49 ( .A1(port0[29]), .A2(n11), .B1(port1[29]), .B2(n13), .ZN(n52)
         );
  AOI22_X1 U50 ( .A1(port0[14]), .A2(n2), .B1(port1[14]), .B2(n12), .ZN(n22)
         );
  AOI22_X1 U51 ( .A1(port0[15]), .A2(n2), .B1(port1[15]), .B2(n14), .ZN(n23)
         );
  AOI22_X1 U52 ( .A1(port0[12]), .A2(n2), .B1(port1[12]), .B2(n15), .ZN(n20)
         );
  AOI22_X1 U53 ( .A1(port0[10]), .A2(n2), .B1(port1[10]), .B2(n12), .ZN(n18)
         );
  AOI22_X1 U54 ( .A1(n1), .A2(port0[27]), .B1(port1[27]), .B2(n15), .ZN(n49)
         );
  AOI22_X1 U55 ( .A1(port0[9]), .A2(n2), .B1(port1[9]), .B2(n12), .ZN(n17) );
  AOI22_X1 U56 ( .A1(port0[24]), .A2(n1), .B1(port1[24]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U57 ( .A1(port0[25]), .A2(n1), .B1(port1[25]), .B2(n15), .ZN(n35)
         );
  AOI22_X1 U58 ( .A1(n11), .A2(port0[0]), .B1(n7), .B2(port1[0]), .ZN(n26) );
  AOI22_X1 U59 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n12), .ZN(n29)
         );
  AOI22_X1 U60 ( .A1(n1), .A2(port0[28]), .B1(port1[28]), .B2(n13), .ZN(n51)
         );
  AOI22_X1 U61 ( .A1(port0[13]), .A2(n3), .B1(port1[13]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U62 ( .A1(port0[22]), .A2(n6), .B1(port1[22]), .B2(n12), .ZN(n31)
         );
  AOI22_X1 U63 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n14), .ZN(n28)
         );
  AOI22_X1 U64 ( .A1(port0[11]), .A2(n6), .B1(port1[11]), .B2(n15), .ZN(n19)
         );
  AOI22_X1 U65 ( .A1(port0[17]), .A2(n6), .B1(port1[17]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U66 ( .A1(port0[16]), .A2(n5), .B1(port1[16]), .B2(n12), .ZN(n24)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n5), .B1(port1[18]), .B2(n12), .ZN(n27)
         );
  AOI22_X1 U68 ( .A1(port0[23]), .A2(n6), .B1(port1[23]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U69 ( .A1(port0[8]), .A2(n6), .B1(port1[8]), .B2(n15), .ZN(n16) );
  INV_X1 U70 ( .A(n56), .ZN(N5) );
  AOI22_X1 U71 ( .A1(port0[5]), .A2(n3), .B1(port1[5]), .B2(n12), .ZN(n58) );
  AOI22_X1 U72 ( .A1(port0[6]), .A2(n5), .B1(port1[6]), .B2(n14), .ZN(n59) );
  AOI22_X1 U73 ( .A1(n4), .A2(port0[30]), .B1(port1[30]), .B2(n13), .ZN(n53)
         );
  AOI22_X1 U74 ( .A1(port0[7]), .A2(n5), .B1(n15), .B2(port1[7]), .ZN(n60) );
  AOI22_X1 U75 ( .A1(port0[2]), .A2(n11), .B1(n13), .B2(port1[2]), .ZN(n55) );
  AOI22_X1 U76 ( .A1(port0[4]), .A2(n6), .B1(port1[4]), .B2(n14), .ZN(n57) );
  AOI22_X1 U77 ( .A1(port0[31]), .A2(n11), .B1(port1[31]), .B2(n8), .ZN(n54)
         );
  AOI22_X1 U78 ( .A1(port0[3]), .A2(n1), .B1(n13), .B2(port1[3]), .ZN(n56) );
  INV_X1 U79 ( .A(n54), .ZN(N33) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_132 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, n41, n45, net140465, net140459, net140457, net140451,
         net140449, net140447, net140495, net169333, net169550, net169651, n1,
         n2, n3, n4, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n35, n38, n39, n40;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  BUF_X1 U1 ( .A(net140495), .Z(net140451) );
  BUF_X1 U2 ( .A(net140451), .Z(n1) );
  BUF_X2 U3 ( .A(sel), .Z(net140495) );
  CLKBUF_X1 U4 ( .A(net140465), .Z(n2) );
  BUF_X1 U5 ( .A(net140495), .Z(net140459) );
  BUF_X2 U6 ( .A(net140495), .Z(net140457) );
  NAND2_X1 U7 ( .A1(port0[3]), .A2(net140449), .ZN(n3) );
  NAND2_X1 U8 ( .A1(port1[3]), .A2(net140451), .ZN(n4) );
  NAND2_X1 U9 ( .A1(n4), .A2(n3), .ZN(portY[3]) );
  CLKBUF_X1 U10 ( .A(sel), .Z(n8) );
  AOI22_X1 U11 ( .A1(n9), .A2(port0[0]), .B1(n7), .B2(port1[0]), .ZN(n6) );
  INV_X1 U12 ( .A(n6), .ZN(N2) );
  BUF_X1 U13 ( .A(n8), .Z(n7) );
  AOI22_X1 U14 ( .A1(port0[1]), .A2(net140447), .B1(net140495), .B2(port1[1]), 
        .ZN(n45) );
  BUF_X1 U15 ( .A(n8), .Z(net140465) );
  INV_X1 U16 ( .A(net140495), .ZN(n9) );
  AOI22_X1 U17 ( .A1(port0[31]), .A2(n9), .B1(port1[31]), .B2(n7), .ZN(n41) );
  INV_X1 U18 ( .A(sel), .ZN(net140447) );
  INV_X1 U19 ( .A(net140457), .ZN(net169651) );
  INV_X1 U20 ( .A(net140457), .ZN(net169550) );
  INV_X1 U21 ( .A(net140451), .ZN(net169333) );
  INV_X1 U22 ( .A(n35), .ZN(N6) );
  INV_X1 U23 ( .A(n33), .ZN(N4) );
  INV_X1 U24 ( .A(n40), .ZN(N9) );
  INV_X1 U25 ( .A(n38), .ZN(N7) );
  INV_X1 U26 ( .A(n24), .ZN(N24) );
  INV_X1 U27 ( .A(n23), .ZN(N23) );
  INV_X1 U28 ( .A(n25), .ZN(N25) );
  INV_X1 U29 ( .A(n17), .ZN(N17) );
  INV_X1 U30 ( .A(n21), .ZN(N21) );
  INV_X1 U31 ( .A(n10), .ZN(N10) );
  INV_X1 U32 ( .A(n14), .ZN(N14) );
  INV_X1 U33 ( .A(n13), .ZN(N13) );
  INV_X1 U34 ( .A(n29), .ZN(N29) );
  INV_X1 U35 ( .A(n27), .ZN(N27) );
  INV_X1 U36 ( .A(n28), .ZN(N28) );
  INV_X1 U37 ( .A(n31), .ZN(N31) );
  INV_X1 U38 ( .A(n16), .ZN(N16) );
  INV_X1 U39 ( .A(n39), .ZN(N8) );
  INV_X1 U40 ( .A(n22), .ZN(N22) );
  INV_X1 U41 ( .A(n30), .ZN(N30) );
  INV_X1 U42 ( .A(n15), .ZN(N15) );
  INV_X1 U43 ( .A(n12), .ZN(N12) );
  INV_X1 U44 ( .A(n11), .ZN(N11) );
  INV_X1 U45 ( .A(n20), .ZN(N20) );
  INV_X1 U46 ( .A(n18), .ZN(N18) );
  INV_X1 U47 ( .A(n19), .ZN(N19) );
  AOI22_X1 U48 ( .A1(port0[26]), .A2(net140447), .B1(port1[26]), .B2(net140451), .ZN(n28) );
  AOI22_X1 U49 ( .A1(port0[22]), .A2(net140447), .B1(port1[22]), .B2(net140457), .ZN(n24) );
  AOI22_X1 U50 ( .A1(port0[21]), .A2(net140447), .B1(port1[21]), .B2(net140457), .ZN(n23) );
  AOI22_X1 U51 ( .A1(port0[29]), .A2(net140447), .B1(net140459), .B2(port1[29]), .ZN(n31) );
  AOI22_X1 U52 ( .A1(port0[23]), .A2(net140447), .B1(port1[23]), .B2(net140457), .ZN(n25) );
  AOI22_X1 U53 ( .A1(port0[20]), .A2(net140447), .B1(port1[20]), .B2(net140451), .ZN(n22) );
  AOI22_X1 U54 ( .A1(port0[28]), .A2(net140447), .B1(net140465), .B2(port1[28]), .ZN(n30) );
  AOI22_X1 U55 ( .A1(port0[19]), .A2(net140447), .B1(port1[19]), .B2(net140457), .ZN(n21) );
  AOI22_X1 U56 ( .A1(port0[27]), .A2(net140447), .B1(net140459), .B2(port1[27]), .ZN(n29) );
  AOI22_X1 U57 ( .A1(port0[25]), .A2(net140447), .B1(port1[25]), .B2(net140451), .ZN(n27) );
  AOI22_X1 U58 ( .A1(port0[24]), .A2(net140447), .B1(port1[24]), .B2(net140457), .ZN(n26) );
  INV_X1 U59 ( .A(n45), .ZN(N3) );
  INV_X1 U60 ( .A(n26), .ZN(N26) );
  INV_X1 U61 ( .A(n32), .ZN(N32) );
  INV_X1 U62 ( .A(net140495), .ZN(net140449) );
  AOI22_X1 U63 ( .A1(port0[13]), .A2(net169550), .B1(port1[13]), .B2(net140457), .ZN(n15) );
  AOI22_X1 U64 ( .A1(port0[17]), .A2(net169333), .B1(port1[17]), .B2(net140457), .ZN(n19) );
  AOI22_X1 U65 ( .A1(port0[12]), .A2(net169651), .B1(port1[12]), .B2(n1), .ZN(
        n14) );
  AOI22_X1 U66 ( .A1(port0[9]), .A2(net169651), .B1(port1[9]), .B2(net140465), 
        .ZN(n11) );
  AOI22_X1 U67 ( .A1(port0[11]), .A2(net169550), .B1(port1[11]), .B2(n1), .ZN(
        n13) );
  AOI22_X1 U68 ( .A1(port0[14]), .A2(net169550), .B1(port1[14]), .B2(n1), .ZN(
        n16) );
  AOI22_X1 U69 ( .A1(port0[10]), .A2(net169651), .B1(port1[10]), .B2(n2), .ZN(
        n12) );
  AOI22_X1 U70 ( .A1(port0[8]), .A2(net169651), .B1(port1[8]), .B2(n2), .ZN(
        n10) );
  AOI22_X1 U71 ( .A1(port0[16]), .A2(net169651), .B1(port1[16]), .B2(net140457), .ZN(n18) );
  AOI22_X1 U72 ( .A1(port0[15]), .A2(net169651), .B1(port1[15]), .B2(n1), .ZN(
        n17) );
  AOI22_X1 U73 ( .A1(port0[18]), .A2(net169550), .B1(port1[18]), .B2(n1), .ZN(
        n20) );
  AOI22_X1 U74 ( .A1(port0[5]), .A2(net169333), .B1(port1[5]), .B2(n2), .ZN(
        n38) );
  AOI22_X1 U75 ( .A1(port0[6]), .A2(net169333), .B1(port1[6]), .B2(net140457), 
        .ZN(n39) );
  AOI22_X1 U76 ( .A1(port0[30]), .A2(net140449), .B1(net140465), .B2(port1[30]), .ZN(n32) );
  AOI22_X1 U77 ( .A1(port0[2]), .A2(net140449), .B1(net140459), .B2(port1[2]), 
        .ZN(n33) );
  AOI22_X1 U78 ( .A1(port0[7]), .A2(net140449), .B1(net140465), .B2(port1[7]), 
        .ZN(n40) );
  AOI22_X1 U79 ( .A1(port0[4]), .A2(net140449), .B1(port1[4]), .B2(net140457), 
        .ZN(n35) );
  INV_X1 U80 ( .A(n41), .ZN(N33) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_131 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16, N17,
         N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30, N31,
         N32, N33, n41, net140435, net140433, net140429, net140427, net140425,
         net140423, net140421, net140419, net140417, net140415, net140439, n1,
         n2, n3, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n35, n37, n38;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  BUF_X1 U1 ( .A(sel), .Z(n1) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n6) );
  BUF_X2 U3 ( .A(net140425), .Z(net140427) );
  BUF_X2 U4 ( .A(sel), .Z(net140439) );
  INV_X1 U5 ( .A(net140439), .ZN(net140419) );
  BUF_X1 U6 ( .A(n1), .Z(net140429) );
  NAND2_X1 U7 ( .A1(port0[0]), .A2(net140417), .ZN(n2) );
  NAND2_X1 U8 ( .A1(port1[0]), .A2(n5), .ZN(n3) );
  NAND2_X1 U9 ( .A1(n2), .A2(n3), .ZN(portY[0]) );
  BUF_X1 U10 ( .A(n1), .Z(net140421) );
  INV_X2 U11 ( .A(net140439), .ZN(net140415) );
  CLKBUF_X1 U12 ( .A(n6), .Z(n5) );
  AOI22_X1 U13 ( .A1(port0[31]), .A2(net140417), .B1(port1[31]), .B2(n5), .ZN(
        n41) );
  BUF_X2 U14 ( .A(n6), .Z(net140425) );
  INV_X1 U15 ( .A(n1), .ZN(net140417) );
  CLKBUF_X1 U16 ( .A(net140439), .Z(net140433) );
  BUF_X2 U17 ( .A(net140439), .Z(net140423) );
  CLKBUF_X1 U18 ( .A(net140433), .Z(net140435) );
  AOI22_X1 U19 ( .A1(port0[24]), .A2(net140419), .B1(port1[24]), .B2(net140427), .ZN(n23) );
  INV_X1 U20 ( .A(n31), .ZN(N4) );
  INV_X1 U21 ( .A(n38), .ZN(N9) );
  INV_X1 U22 ( .A(n35), .ZN(N7) );
  INV_X1 U23 ( .A(n21), .ZN(N24) );
  AOI22_X1 U24 ( .A1(port0[22]), .A2(net140419), .B1(port1[22]), .B2(net140427), .ZN(n21) );
  INV_X1 U25 ( .A(n20), .ZN(N23) );
  AOI22_X1 U26 ( .A1(port0[21]), .A2(net140415), .B1(port1[21]), .B2(net140427), .ZN(n20) );
  INV_X1 U27 ( .A(n22), .ZN(N25) );
  AOI22_X1 U28 ( .A1(port0[23]), .A2(net140415), .B1(port1[23]), .B2(net140427), .ZN(n22) );
  INV_X1 U29 ( .A(n14), .ZN(N17) );
  AOI22_X1 U30 ( .A1(port0[15]), .A2(net140415), .B1(port1[15]), .B2(net140423), .ZN(n14) );
  INV_X1 U31 ( .A(n18), .ZN(N21) );
  AOI22_X1 U32 ( .A1(port0[19]), .A2(net140415), .B1(port1[19]), .B2(net140429), .ZN(n18) );
  INV_X1 U33 ( .A(n7), .ZN(N10) );
  AOI22_X1 U34 ( .A1(port0[8]), .A2(net140415), .B1(port1[8]), .B2(net140435), 
        .ZN(n7) );
  INV_X1 U35 ( .A(n11), .ZN(N14) );
  AOI22_X1 U36 ( .A1(port0[12]), .A2(net140415), .B1(port1[12]), .B2(net140433), .ZN(n11) );
  INV_X1 U37 ( .A(n10), .ZN(N13) );
  AOI22_X1 U38 ( .A1(port0[11]), .A2(net140415), .B1(port1[11]), .B2(net140433), .ZN(n10) );
  INV_X1 U39 ( .A(n26), .ZN(N29) );
  AOI22_X1 U40 ( .A1(port0[27]), .A2(net140419), .B1(port1[27]), .B2(net140425), .ZN(n26) );
  INV_X1 U41 ( .A(n24), .ZN(N27) );
  AOI22_X1 U42 ( .A1(port0[25]), .A2(net140419), .B1(port1[25]), .B2(net140425), .ZN(n24) );
  INV_X1 U43 ( .A(n25), .ZN(N28) );
  INV_X1 U44 ( .A(n29), .ZN(N31) );
  INV_X1 U45 ( .A(n13), .ZN(N16) );
  INV_X1 U46 ( .A(n37), .ZN(N8) );
  INV_X1 U47 ( .A(n19), .ZN(N22) );
  INV_X1 U48 ( .A(n28), .ZN(N30) );
  INV_X1 U49 ( .A(n12), .ZN(N15) );
  INV_X1 U50 ( .A(n9), .ZN(N12) );
  INV_X1 U51 ( .A(n8), .ZN(N11) );
  INV_X1 U52 ( .A(n17), .ZN(N20) );
  INV_X1 U53 ( .A(n15), .ZN(N18) );
  INV_X1 U54 ( .A(n16), .ZN(N19) );
  AOI22_X1 U55 ( .A1(port0[20]), .A2(net140415), .B1(port1[20]), .B2(net140429), .ZN(n19) );
  AOI22_X1 U56 ( .A1(port0[13]), .A2(net140415), .B1(port1[13]), .B2(net140433), .ZN(n12) );
  AOI22_X1 U57 ( .A1(port0[26]), .A2(net140415), .B1(port1[26]), .B2(net140425), .ZN(n25) );
  AOI22_X1 U58 ( .A1(port0[28]), .A2(net140419), .B1(port1[28]), .B2(net140423), .ZN(n28) );
  AOI22_X1 U59 ( .A1(port0[10]), .A2(net140415), .B1(port1[10]), .B2(net140435), .ZN(n9) );
  AOI22_X1 U60 ( .A1(port0[17]), .A2(net140415), .B1(port1[17]), .B2(net140423), .ZN(n16) );
  AOI22_X1 U61 ( .A1(port0[16]), .A2(net140415), .B1(port1[16]), .B2(net140423), .ZN(n15) );
  AOI22_X1 U62 ( .A1(port0[14]), .A2(net140415), .B1(port1[14]), .B2(net140433), .ZN(n13) );
  AOI22_X1 U63 ( .A1(port0[18]), .A2(net140415), .B1(port1[18]), .B2(net140429), .ZN(n17) );
  AOI22_X1 U64 ( .A1(port0[9]), .A2(net140415), .B1(port1[9]), .B2(net140435), 
        .ZN(n8) );
  AOI22_X1 U65 ( .A1(port0[29]), .A2(net140419), .B1(port1[29]), .B2(net140429), .ZN(n29) );
  AOI22_X1 U66 ( .A1(port0[1]), .A2(net140417), .B1(port1[1]), .B2(net140425), 
        .ZN(n27) );
  INV_X1 U67 ( .A(n27), .ZN(N3) );
  INV_X1 U68 ( .A(n33), .ZN(N6) );
  INV_X1 U69 ( .A(n23), .ZN(N26) );
  AOI22_X1 U70 ( .A1(port0[30]), .A2(net140417), .B1(port1[30]), .B2(net140423), .ZN(n30) );
  AOI22_X1 U71 ( .A1(port0[2]), .A2(net140419), .B1(port1[2]), .B2(net140423), 
        .ZN(n31) );
  AOI22_X1 U72 ( .A1(port0[5]), .A2(net140415), .B1(port1[5]), .B2(net140421), 
        .ZN(n35) );
  AOI22_X1 U73 ( .A1(port0[6]), .A2(net140415), .B1(port1[6]), .B2(net140421), 
        .ZN(n37) );
  AOI22_X1 U74 ( .A1(port0[7]), .A2(net140415), .B1(net140435), .B2(port1[7]), 
        .ZN(n38) );
  AOI22_X1 U75 ( .A1(port0[4]), .A2(net140415), .B1(port1[4]), .B2(net140421), 
        .ZN(n33) );
  INV_X1 U76 ( .A(n30), .ZN(N32) );
  INV_X1 U77 ( .A(n32), .ZN(N5) );
  AOI22_X1 U78 ( .A1(port0[3]), .A2(net140419), .B1(port1[3]), .B2(net140421), 
        .ZN(n32) );
  INV_X1 U79 ( .A(n41), .ZN(N33) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_130 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, n57, n58, n59, net132559, net132557, net132553, net132551,
         net132549, net132547, net132545, net132543, net132541, net132539,
         net132579, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;

  MUX2_X2 U1 ( .A(port0[1]), .B(port1[1]), .S(sel), .Z(N3) );
  MUX2_X2 U2 ( .A(port1[0]), .B(port0[0]), .S(net132543), .Z(N2) );
  INV_X2 U3 ( .A(n5), .ZN(net132543) );
  NAND2_X1 U4 ( .A1(port0[31]), .A2(net132543), .ZN(n1) );
  NAND2_X1 U5 ( .A1(port1[31]), .A2(net132547), .ZN(n2) );
  NAND2_X1 U6 ( .A1(n2), .A2(n1), .ZN(portY[31]) );
  BUF_X1 U7 ( .A(n6), .Z(n4) );
  AOI22_X1 U8 ( .A1(port0[15]), .A2(net132539), .B1(port1[15]), .B2(n4), .ZN(
        n59) );
  AOI22_X1 U9 ( .A1(port0[17]), .A2(net132539), .B1(port1[17]), .B2(n4), .ZN(
        n57) );
  AOI22_X1 U10 ( .A1(port0[16]), .A2(net132539), .B1(port1[16]), .B2(n4), .ZN(
        n58) );
  CLKBUF_X1 U11 ( .A(sel), .Z(n6) );
  BUF_X1 U12 ( .A(n6), .Z(net132551) );
  BUF_X1 U13 ( .A(n6), .Z(net132553) );
  INV_X1 U14 ( .A(n5), .ZN(net132539) );
  BUF_X1 U15 ( .A(n7), .Z(n5) );
  INV_X1 U16 ( .A(n5), .ZN(net132541) );
  CLKBUF_X1 U17 ( .A(sel), .Z(n7) );
  CLKBUF_X1 U18 ( .A(n7), .Z(net132557) );
  CLKBUF_X1 U19 ( .A(n7), .Z(net132559) );
  CLKBUF_X1 U20 ( .A(sel), .Z(net132579) );
  BUF_X1 U21 ( .A(net132579), .Z(net132547) );
  AOI22_X1 U22 ( .A1(port0[30]), .A2(net132543), .B1(port1[30]), .B2(net132547), .ZN(n27) );
  AOI22_X1 U23 ( .A1(port0[24]), .A2(net132541), .B1(port1[24]), .B2(net132551), .ZN(n21) );
  INV_X1 U24 ( .A(n29), .ZN(N5) );
  INV_X1 U25 ( .A(n30), .ZN(N6) );
  INV_X1 U26 ( .A(n33), .ZN(N9) );
  AOI22_X1 U27 ( .A1(port0[7]), .A2(net132543), .B1(net132559), .B2(port1[7]), 
        .ZN(n33) );
  INV_X1 U28 ( .A(n28), .ZN(N4) );
  AOI22_X1 U29 ( .A1(port0[2]), .A2(net132543), .B1(port1[2]), .B2(net132547), 
        .ZN(n28) );
  INV_X1 U30 ( .A(n31), .ZN(N7) );
  AOI22_X1 U31 ( .A1(port0[5]), .A2(net132543), .B1(port1[5]), .B2(net132545), 
        .ZN(n31) );
  INV_X1 U32 ( .A(n32), .ZN(N8) );
  AOI22_X1 U33 ( .A1(port0[6]), .A2(net132543), .B1(port1[6]), .B2(net132545), 
        .ZN(n32) );
  INV_X1 U34 ( .A(n9), .ZN(N11) );
  AOI22_X1 U35 ( .A1(port0[9]), .A2(net132539), .B1(port1[9]), .B2(net132559), 
        .ZN(n9) );
  INV_X1 U36 ( .A(n59), .ZN(N17) );
  INV_X1 U37 ( .A(n19), .ZN(N24) );
  AOI22_X1 U38 ( .A1(port0[22]), .A2(net132541), .B1(port1[22]), .B2(net132551), .ZN(n19) );
  INV_X1 U39 ( .A(n8), .ZN(N10) );
  AOI22_X1 U40 ( .A1(port0[8]), .A2(net132539), .B1(port1[8]), .B2(net132559), 
        .ZN(n8) );
  INV_X1 U41 ( .A(n11), .ZN(N13) );
  AOI22_X1 U42 ( .A1(port0[11]), .A2(net132539), .B1(port1[11]), .B2(net132557), .ZN(n11) );
  INV_X1 U43 ( .A(n20), .ZN(N25) );
  AOI22_X1 U44 ( .A1(port0[23]), .A2(net132541), .B1(port1[23]), .B2(net132551), .ZN(n20) );
  INV_X1 U45 ( .A(n12), .ZN(N14) );
  AOI22_X1 U46 ( .A1(port0[12]), .A2(net132539), .B1(port1[12]), .B2(net132557), .ZN(n12) );
  INV_X1 U47 ( .A(n22), .ZN(N27) );
  AOI22_X1 U48 ( .A1(port0[25]), .A2(net132541), .B1(port1[25]), .B2(net132549), .ZN(n22) );
  INV_X1 U49 ( .A(n16), .ZN(N21) );
  AOI22_X1 U50 ( .A1(port0[19]), .A2(net132541), .B1(port1[19]), .B2(net132553), .ZN(n16) );
  INV_X1 U51 ( .A(n18), .ZN(N23) );
  AOI22_X1 U52 ( .A1(port0[21]), .A2(net132541), .B1(port1[21]), .B2(net132551), .ZN(n18) );
  INV_X1 U53 ( .A(n24), .ZN(N29) );
  AOI22_X1 U54 ( .A1(port0[27]), .A2(net132541), .B1(port1[27]), .B2(net132549), .ZN(n24) );
  INV_X1 U55 ( .A(n10), .ZN(N12) );
  AOI22_X1 U56 ( .A1(port0[10]), .A2(net132539), .B1(port1[10]), .B2(net132559), .ZN(n10) );
  INV_X1 U57 ( .A(n57), .ZN(N19) );
  INV_X1 U58 ( .A(n15), .ZN(N20) );
  AOI22_X1 U59 ( .A1(port0[18]), .A2(net132539), .B1(port1[18]), .B2(net132553), .ZN(n15) );
  INV_X1 U60 ( .A(n58), .ZN(N18) );
  INV_X1 U61 ( .A(n13), .ZN(N15) );
  AOI22_X1 U62 ( .A1(port0[13]), .A2(net132539), .B1(port1[13]), .B2(net132557), .ZN(n13) );
  INV_X1 U63 ( .A(n14), .ZN(N16) );
  AOI22_X1 U64 ( .A1(port0[14]), .A2(net132539), .B1(port1[14]), .B2(net132557), .ZN(n14) );
  INV_X1 U65 ( .A(n25), .ZN(N30) );
  AOI22_X1 U66 ( .A1(port0[28]), .A2(net132541), .B1(port1[28]), .B2(net132547), .ZN(n25) );
  INV_X1 U67 ( .A(n17), .ZN(N22) );
  AOI22_X1 U68 ( .A1(port0[20]), .A2(net132541), .B1(port1[20]), .B2(net132553), .ZN(n17) );
  INV_X1 U69 ( .A(n26), .ZN(N31) );
  AOI22_X1 U70 ( .A1(port0[29]), .A2(net132541), .B1(port1[29]), .B2(net132553), .ZN(n26) );
  INV_X1 U71 ( .A(n23), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(net132541), .B1(port1[26]), .B2(net132549), .ZN(n23) );
  CLKBUF_X1 U73 ( .A(net132579), .Z(net132549) );
  CLKBUF_X1 U74 ( .A(net132579), .Z(net132545) );
  AOI22_X1 U75 ( .A1(port0[4]), .A2(net132543), .B1(port1[4]), .B2(net132545), 
        .ZN(n30) );
  INV_X1 U76 ( .A(n21), .ZN(N26) );
  INV_X1 U77 ( .A(n27), .ZN(N32) );
  AOI22_X1 U78 ( .A1(port0[3]), .A2(net132543), .B1(port1[3]), .B2(net132545), 
        .ZN(n29) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_129 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N28, N30, N32, N33,
         n1, n2, n4, n5, n7, n8, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32,
         n33, n35, n41, n43, n46, n48, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[26] = N28;
  assign portY[28] = N30;
  assign portY[30] = N32;
  assign portY[31] = N33;

  MUX2_X1 U1 ( .A(port0[31]), .B(port1[31]), .S(sel), .Z(N33) );
  NAND2_X1 U2 ( .A1(port0[25]), .A2(n14), .ZN(n1) );
  NAND2_X1 U3 ( .A1(port1[25]), .A2(n18), .ZN(n2) );
  NAND2_X1 U4 ( .A1(n1), .A2(n2), .ZN(portY[25]) );
  NAND2_X1 U5 ( .A1(port0[27]), .A2(n14), .ZN(n4) );
  NAND2_X1 U6 ( .A1(port1[27]), .A2(n18), .ZN(n5) );
  NAND2_X1 U7 ( .A1(n4), .A2(n5), .ZN(portY[27]) );
  INV_X2 U8 ( .A(n24), .ZN(n14) );
  NAND2_X1 U9 ( .A1(port0[29]), .A2(n14), .ZN(n7) );
  NAND2_X1 U10 ( .A1(port1[29]), .A2(n20), .ZN(n8) );
  NAND2_X1 U11 ( .A1(n7), .A2(n8), .ZN(portY[29]) );
  CLKBUF_X1 U12 ( .A(n12), .Z(n22) );
  CLKBUF_X1 U13 ( .A(n11), .Z(n19) );
  CLKBUF_X1 U14 ( .A(n10), .Z(n18) );
  BUF_X1 U15 ( .A(n12), .Z(n24) );
  INV_X1 U16 ( .A(n24), .ZN(n13) );
  INV_X1 U17 ( .A(n66), .ZN(N9) );
  AOI22_X1 U18 ( .A1(port0[7]), .A2(n15), .B1(n23), .B2(port1[7]), .ZN(n66) );
  INV_X1 U19 ( .A(n33), .ZN(N18) );
  AOI22_X1 U20 ( .A1(port0[16]), .A2(n13), .B1(port1[16]), .B2(n21), .ZN(n33)
         );
  INV_X1 U21 ( .A(n35), .ZN(N19) );
  AOI22_X1 U22 ( .A1(port0[17]), .A2(n13), .B1(port1[17]), .B2(n21), .ZN(n35)
         );
  INV_X1 U23 ( .A(n63), .ZN(N6) );
  INV_X1 U24 ( .A(n62), .ZN(N5) );
  INV_X1 U25 ( .A(n64), .ZN(N7) );
  AOI22_X1 U26 ( .A1(port0[5]), .A2(n15), .B1(port1[5]), .B2(n16), .ZN(n64) );
  INV_X1 U27 ( .A(n65), .ZN(N8) );
  AOI22_X1 U28 ( .A1(port0[6]), .A2(n15), .B1(port1[6]), .B2(n16), .ZN(n65) );
  INV_X1 U29 ( .A(n61), .ZN(N4) );
  AOI22_X1 U30 ( .A1(port0[2]), .A2(n15), .B1(port1[2]), .B2(n17), .ZN(n61) );
  INV_X1 U31 ( .A(n26), .ZN(N11) );
  AOI22_X1 U32 ( .A1(port0[9]), .A2(n13), .B1(port1[9]), .B2(n23), .ZN(n26) );
  INV_X1 U33 ( .A(n58), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n14), .B1(port1[1]), .B2(n18), .ZN(n58) );
  INV_X1 U35 ( .A(n54), .ZN(N24) );
  AOI22_X1 U36 ( .A1(port0[22]), .A2(n14), .B1(port1[22]), .B2(n19), .ZN(n54)
         );
  INV_X1 U37 ( .A(n55), .ZN(N25) );
  AOI22_X1 U38 ( .A1(port0[23]), .A2(n14), .B1(port1[23]), .B2(n19), .ZN(n55)
         );
  INV_X1 U39 ( .A(n46), .ZN(N21) );
  AOI22_X1 U40 ( .A1(port0[19]), .A2(n14), .B1(port1[19]), .B2(n20), .ZN(n46)
         );
  INV_X1 U41 ( .A(n29), .ZN(N14) );
  AOI22_X1 U42 ( .A1(port0[12]), .A2(n13), .B1(port1[12]), .B2(n22), .ZN(n29)
         );
  INV_X1 U43 ( .A(n25), .ZN(N10) );
  AOI22_X1 U44 ( .A1(port0[8]), .A2(n13), .B1(port1[8]), .B2(n23), .ZN(n25) );
  INV_X1 U45 ( .A(n28), .ZN(N13) );
  AOI22_X1 U46 ( .A1(port0[11]), .A2(n13), .B1(port1[11]), .B2(n22), .ZN(n28)
         );
  INV_X1 U47 ( .A(n56), .ZN(N26) );
  AOI22_X1 U48 ( .A1(port0[24]), .A2(n14), .B1(port1[24]), .B2(n19), .ZN(n56)
         );
  INV_X1 U49 ( .A(n43), .ZN(N20) );
  AOI22_X1 U50 ( .A1(port0[18]), .A2(n13), .B1(port1[18]), .B2(n20), .ZN(n43)
         );
  INV_X1 U51 ( .A(n57), .ZN(N28) );
  AOI22_X1 U52 ( .A1(port0[26]), .A2(n14), .B1(port1[26]), .B2(n18), .ZN(n57)
         );
  INV_X1 U53 ( .A(n53), .ZN(N23) );
  AOI22_X1 U54 ( .A1(port0[21]), .A2(n14), .B1(port1[21]), .B2(n19), .ZN(n53)
         );
  INV_X1 U55 ( .A(n48), .ZN(N22) );
  AOI22_X1 U56 ( .A1(port0[20]), .A2(n14), .B1(port1[20]), .B2(n20), .ZN(n48)
         );
  INV_X1 U57 ( .A(n59), .ZN(N30) );
  AOI22_X1 U58 ( .A1(port0[28]), .A2(n14), .B1(port1[28]), .B2(n17), .ZN(n59)
         );
  INV_X1 U59 ( .A(n31), .ZN(N16) );
  AOI22_X1 U60 ( .A1(port0[14]), .A2(n13), .B1(port1[14]), .B2(n22), .ZN(n31)
         );
  INV_X1 U61 ( .A(n30), .ZN(N15) );
  AOI22_X1 U62 ( .A1(port0[13]), .A2(n13), .B1(port1[13]), .B2(n22), .ZN(n30)
         );
  INV_X1 U63 ( .A(n32), .ZN(N17) );
  AOI22_X1 U64 ( .A1(port0[15]), .A2(n13), .B1(port1[15]), .B2(n21), .ZN(n32)
         );
  INV_X1 U65 ( .A(n27), .ZN(N12) );
  AOI22_X1 U66 ( .A1(port0[10]), .A2(n13), .B1(port1[10]), .B2(n23), .ZN(n27)
         );
  INV_X1 U67 ( .A(n41), .ZN(N2) );
  AOI22_X1 U68 ( .A1(port0[0]), .A2(n13), .B1(port1[0]), .B2(n21), .ZN(n41) );
  BUF_X1 U69 ( .A(n11), .Z(n20) );
  CLKBUF_X1 U70 ( .A(n11), .Z(n21) );
  CLKBUF_X1 U71 ( .A(n12), .Z(n23) );
  BUF_X1 U72 ( .A(n10), .Z(n17) );
  CLKBUF_X1 U73 ( .A(n10), .Z(n16) );
  CLKBUF_X1 U74 ( .A(sel), .Z(n12) );
  CLKBUF_X1 U75 ( .A(sel), .Z(n10) );
  CLKBUF_X1 U76 ( .A(sel), .Z(n11) );
  AOI22_X1 U77 ( .A1(port0[4]), .A2(n15), .B1(port1[4]), .B2(n16), .ZN(n63) );
  INV_X1 U78 ( .A(n60), .ZN(N32) );
  AOI22_X1 U79 ( .A1(port0[30]), .A2(n15), .B1(port1[30]), .B2(n17), .ZN(n60)
         );
  AOI22_X1 U80 ( .A1(port0[3]), .A2(n15), .B1(port1[3]), .B2(n16), .ZN(n62) );
  INV_X1 U81 ( .A(n24), .ZN(n15) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_128 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  BUF_X1 U3 ( .A(n1), .Z(n6) );
  BUF_X1 U4 ( .A(n3), .Z(n12) );
  BUF_X1 U5 ( .A(n2), .Z(n11) );
  BUF_X1 U6 ( .A(n2), .Z(n9) );
  BUF_X1 U7 ( .A(n1), .Z(n8) );
  BUF_X1 U8 ( .A(n2), .Z(n10) );
  BUF_X1 U9 ( .A(n3), .Z(n14) );
  BUF_X1 U10 ( .A(n3), .Z(n13) );
  BUF_X1 U11 ( .A(n1), .Z(n7) );
  INV_X1 U12 ( .A(n51), .ZN(N32) );
  INV_X1 U13 ( .A(n52), .ZN(N33) );
  BUF_X1 U14 ( .A(sel), .Z(n3) );
  BUF_X1 U15 ( .A(sel), .Z(n2) );
  BUF_X1 U16 ( .A(sel), .Z(n1) );
  INV_X1 U17 ( .A(n23), .ZN(N18) );
  INV_X1 U18 ( .A(n24), .ZN(N19) );
  INV_X1 U19 ( .A(n26), .ZN(N20) );
  INV_X1 U20 ( .A(n27), .ZN(N21) );
  INV_X1 U21 ( .A(n28), .ZN(N22) );
  INV_X1 U22 ( .A(n29), .ZN(N23) );
  INV_X1 U23 ( .A(n30), .ZN(N24) );
  INV_X1 U24 ( .A(n31), .ZN(N25) );
  INV_X1 U25 ( .A(n32), .ZN(N26) );
  INV_X1 U26 ( .A(n33), .ZN(N27) );
  INV_X1 U27 ( .A(n35), .ZN(N28) );
  INV_X1 U28 ( .A(n47), .ZN(N29) );
  INV_X1 U29 ( .A(n49), .ZN(N30) );
  INV_X1 U30 ( .A(n50), .ZN(N31) );
  INV_X1 U31 ( .A(n53), .ZN(N4) );
  AOI22_X1 U32 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U33 ( .A(n54), .ZN(N5) );
  AOI22_X1 U34 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U35 ( .A(n55), .ZN(N6) );
  AOI22_X1 U36 ( .A1(port0[4]), .A2(n5), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U37 ( .A(n56), .ZN(N7) );
  AOI22_X1 U38 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U39 ( .A(n57), .ZN(N8) );
  AOI22_X1 U40 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n6), .ZN(n57) );
  AOI22_X1 U41 ( .A1(port0[30]), .A2(n4), .B1(port1[30]), .B2(n7), .ZN(n51) );
  INV_X1 U42 ( .A(n25), .ZN(N2) );
  AOI22_X1 U43 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  INV_X1 U44 ( .A(n48), .ZN(N3) );
  AOI22_X1 U45 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  AOI22_X1 U46 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  AOI22_X1 U47 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  AOI22_X1 U48 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  AOI22_X1 U49 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  AOI22_X1 U50 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  AOI22_X1 U51 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  AOI22_X1 U52 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  AOI22_X1 U53 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  AOI22_X1 U54 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  AOI22_X1 U55 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  AOI22_X1 U56 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  AOI22_X1 U57 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  AOI22_X1 U58 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  AOI22_X1 U59 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  INV_X1 U60 ( .A(n58), .ZN(N9) );
  AOI22_X1 U61 ( .A1(port0[7]), .A2(n4), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U62 ( .A(n15), .ZN(N10) );
  AOI22_X1 U63 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U64 ( .A(n16), .ZN(N11) );
  AOI22_X1 U65 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U66 ( .A(n17), .ZN(N12) );
  AOI22_X1 U67 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U68 ( .A(n18), .ZN(N13) );
  AOI22_X1 U69 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U70 ( .A(n19), .ZN(N14) );
  AOI22_X1 U71 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U72 ( .A(n20), .ZN(N15) );
  AOI22_X1 U73 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U74 ( .A(n21), .ZN(N16) );
  AOI22_X1 U75 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U76 ( .A(n22), .ZN(N17) );
  AOI22_X1 U77 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  AOI22_X1 U78 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n7), .ZN(n52) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_126 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  BUF_X1 U3 ( .A(n1), .Z(n6) );
  BUF_X1 U4 ( .A(n3), .Z(n12) );
  BUF_X1 U5 ( .A(n2), .Z(n11) );
  BUF_X1 U6 ( .A(n2), .Z(n9) );
  BUF_X1 U7 ( .A(n1), .Z(n8) );
  BUF_X1 U8 ( .A(n2), .Z(n10) );
  BUF_X1 U9 ( .A(n1), .Z(n7) );
  BUF_X1 U10 ( .A(n3), .Z(n14) );
  BUF_X1 U11 ( .A(n3), .Z(n13) );
  BUF_X1 U12 ( .A(sel), .Z(n3) );
  BUF_X1 U13 ( .A(sel), .Z(n2) );
  BUF_X1 U14 ( .A(sel), .Z(n1) );
  INV_X1 U15 ( .A(n53), .ZN(N4) );
  AOI22_X1 U16 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U17 ( .A(n54), .ZN(N5) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U19 ( .A(n55), .ZN(N6) );
  AOI22_X1 U20 ( .A1(port0[4]), .A2(n5), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U21 ( .A(n56), .ZN(N7) );
  AOI22_X1 U22 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U23 ( .A(n57), .ZN(N8) );
  AOI22_X1 U24 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U25 ( .A(n58), .ZN(N9) );
  AOI22_X1 U26 ( .A1(port0[7]), .A2(n4), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U27 ( .A(n51), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n4), .B1(port1[30]), .B2(n7), .ZN(n51) );
  INV_X1 U29 ( .A(n52), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n7), .ZN(n52) );
  INV_X1 U31 ( .A(n25), .ZN(N2) );
  AOI22_X1 U32 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  INV_X1 U33 ( .A(n48), .ZN(N3) );
  AOI22_X1 U34 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  INV_X1 U35 ( .A(n15), .ZN(N10) );
  AOI22_X1 U36 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U37 ( .A(n16), .ZN(N11) );
  AOI22_X1 U38 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U39 ( .A(n17), .ZN(N12) );
  AOI22_X1 U40 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U41 ( .A(n18), .ZN(N13) );
  AOI22_X1 U42 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U43 ( .A(n19), .ZN(N14) );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U45 ( .A(n20), .ZN(N15) );
  AOI22_X1 U46 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U47 ( .A(n21), .ZN(N16) );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U49 ( .A(n22), .ZN(N17) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  INV_X1 U51 ( .A(n23), .ZN(N18) );
  AOI22_X1 U52 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  INV_X1 U53 ( .A(n24), .ZN(N19) );
  AOI22_X1 U54 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U55 ( .A(n26), .ZN(N20) );
  AOI22_X1 U56 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  INV_X1 U57 ( .A(n27), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  INV_X1 U59 ( .A(n28), .ZN(N22) );
  AOI22_X1 U60 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U61 ( .A(n29), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  INV_X1 U63 ( .A(n30), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  INV_X1 U65 ( .A(n31), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  INV_X1 U67 ( .A(n32), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U69 ( .A(n33), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  INV_X1 U71 ( .A(n35), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  INV_X1 U73 ( .A(n47), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  INV_X1 U75 ( .A(n49), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U77 ( .A(n50), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_125 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  BUF_X1 U3 ( .A(n1), .Z(n6) );
  BUF_X1 U4 ( .A(n3), .Z(n12) );
  BUF_X1 U5 ( .A(n2), .Z(n11) );
  BUF_X1 U6 ( .A(n2), .Z(n9) );
  BUF_X1 U7 ( .A(n1), .Z(n8) );
  BUF_X1 U8 ( .A(n2), .Z(n10) );
  BUF_X1 U9 ( .A(n1), .Z(n7) );
  BUF_X1 U10 ( .A(n3), .Z(n14) );
  BUF_X1 U11 ( .A(n3), .Z(n13) );
  BUF_X1 U12 ( .A(sel), .Z(n3) );
  BUF_X1 U13 ( .A(sel), .Z(n2) );
  BUF_X1 U14 ( .A(sel), .Z(n1) );
  INV_X1 U15 ( .A(n52), .ZN(N33) );
  AOI22_X1 U16 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n7), .ZN(n52) );
  INV_X1 U17 ( .A(n51), .ZN(N32) );
  AOI22_X1 U18 ( .A1(port0[30]), .A2(n4), .B1(port1[30]), .B2(n7), .ZN(n51) );
  INV_X1 U19 ( .A(n50), .ZN(N31) );
  AOI22_X1 U20 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  INV_X1 U21 ( .A(n49), .ZN(N30) );
  AOI22_X1 U22 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U23 ( .A(n47), .ZN(N29) );
  AOI22_X1 U24 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  INV_X1 U25 ( .A(n35), .ZN(N28) );
  AOI22_X1 U26 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  INV_X1 U27 ( .A(n58), .ZN(N9) );
  AOI22_X1 U28 ( .A1(port0[7]), .A2(n4), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U29 ( .A(n33), .ZN(N27) );
  AOI22_X1 U30 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  INV_X1 U31 ( .A(n32), .ZN(N26) );
  AOI22_X1 U32 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U33 ( .A(n31), .ZN(N25) );
  AOI22_X1 U34 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  INV_X1 U35 ( .A(n30), .ZN(N24) );
  AOI22_X1 U36 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  INV_X1 U37 ( .A(n29), .ZN(N23) );
  AOI22_X1 U38 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  INV_X1 U39 ( .A(n28), .ZN(N22) );
  AOI22_X1 U40 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U41 ( .A(n27), .ZN(N21) );
  AOI22_X1 U42 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  INV_X1 U43 ( .A(n26), .ZN(N20) );
  AOI22_X1 U44 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  INV_X1 U45 ( .A(n20), .ZN(N15) );
  AOI22_X1 U46 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U47 ( .A(n21), .ZN(N16) );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U49 ( .A(n24), .ZN(N19) );
  AOI22_X1 U50 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U51 ( .A(n23), .ZN(N18) );
  AOI22_X1 U52 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  INV_X1 U53 ( .A(n22), .ZN(N17) );
  AOI22_X1 U54 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  INV_X1 U55 ( .A(n55), .ZN(N6) );
  AOI22_X1 U56 ( .A1(port0[4]), .A2(n5), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U57 ( .A(n56), .ZN(N7) );
  AOI22_X1 U58 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U59 ( .A(n57), .ZN(N8) );
  AOI22_X1 U60 ( .A1(port0[6]), .A2(n5), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U61 ( .A(n15), .ZN(N10) );
  AOI22_X1 U62 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U63 ( .A(n16), .ZN(N11) );
  AOI22_X1 U64 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U65 ( .A(n17), .ZN(N12) );
  AOI22_X1 U66 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U67 ( .A(n18), .ZN(N13) );
  AOI22_X1 U68 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U69 ( .A(n19), .ZN(N14) );
  AOI22_X1 U70 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U71 ( .A(n48), .ZN(N3) );
  AOI22_X1 U72 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  INV_X1 U73 ( .A(n53), .ZN(N4) );
  AOI22_X1 U74 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U75 ( .A(n54), .ZN(N5) );
  AOI22_X1 U76 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U77 ( .A(n25), .ZN(N2) );
  AOI22_X1 U78 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_124 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n5) );
  INV_X1 U2 ( .A(n14), .ZN(n4) );
  BUF_X1 U3 ( .A(n2), .Z(n9) );
  BUF_X1 U4 ( .A(n2), .Z(n10) );
  BUF_X1 U5 ( .A(n3), .Z(n12) );
  BUF_X1 U6 ( .A(n1), .Z(n6) );
  BUF_X1 U7 ( .A(n1), .Z(n7) );
  BUF_X1 U8 ( .A(n1), .Z(n8) );
  BUF_X1 U9 ( .A(n2), .Z(n11) );
  BUF_X1 U10 ( .A(n3), .Z(n14) );
  BUF_X1 U11 ( .A(n3), .Z(n13) );
  BUF_X1 U12 ( .A(sel), .Z(n3) );
  BUF_X1 U13 ( .A(sel), .Z(n1) );
  BUF_X1 U14 ( .A(sel), .Z(n2) );
  INV_X1 U15 ( .A(n52), .ZN(N33) );
  AOI22_X1 U16 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n7), .ZN(n52) );
  INV_X1 U17 ( .A(n51), .ZN(N32) );
  AOI22_X1 U18 ( .A1(port0[30]), .A2(n4), .B1(port1[30]), .B2(n7), .ZN(n51) );
  INV_X1 U19 ( .A(n50), .ZN(N31) );
  AOI22_X1 U20 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  INV_X1 U21 ( .A(n49), .ZN(N30) );
  AOI22_X1 U22 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U23 ( .A(n47), .ZN(N29) );
  AOI22_X1 U24 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  INV_X1 U25 ( .A(n35), .ZN(N28) );
  AOI22_X1 U26 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  INV_X1 U27 ( .A(n33), .ZN(N27) );
  AOI22_X1 U28 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  INV_X1 U29 ( .A(n32), .ZN(N26) );
  AOI22_X1 U30 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U31 ( .A(n31), .ZN(N25) );
  AOI22_X1 U32 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  INV_X1 U33 ( .A(n30), .ZN(N24) );
  AOI22_X1 U34 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  INV_X1 U35 ( .A(n29), .ZN(N23) );
  AOI22_X1 U36 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  INV_X1 U37 ( .A(n28), .ZN(N22) );
  AOI22_X1 U38 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U39 ( .A(n27), .ZN(N21) );
  AOI22_X1 U40 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  INV_X1 U41 ( .A(n26), .ZN(N20) );
  AOI22_X1 U42 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  INV_X1 U43 ( .A(n24), .ZN(N19) );
  AOI22_X1 U44 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U45 ( .A(n23), .ZN(N18) );
  AOI22_X1 U46 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  INV_X1 U47 ( .A(n22), .ZN(N17) );
  AOI22_X1 U48 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  INV_X1 U49 ( .A(n21), .ZN(N16) );
  AOI22_X1 U50 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U51 ( .A(n20), .ZN(N15) );
  AOI22_X1 U52 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U53 ( .A(n19), .ZN(N14) );
  AOI22_X1 U54 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U55 ( .A(n18), .ZN(N13) );
  AOI22_X1 U56 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U57 ( .A(n17), .ZN(N12) );
  AOI22_X1 U58 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U59 ( .A(n16), .ZN(N11) );
  AOI22_X1 U60 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U61 ( .A(n15), .ZN(N10) );
  AOI22_X1 U62 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U63 ( .A(n58), .ZN(N9) );
  AOI22_X1 U64 ( .A1(port0[7]), .A2(n4), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U65 ( .A(n57), .ZN(N8) );
  AOI22_X1 U66 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U67 ( .A(n56), .ZN(N7) );
  AOI22_X1 U68 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U69 ( .A(n55), .ZN(N6) );
  AOI22_X1 U70 ( .A1(port0[4]), .A2(n5), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U71 ( .A(n54), .ZN(N5) );
  AOI22_X1 U72 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U73 ( .A(n53), .ZN(N4) );
  AOI22_X1 U74 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U75 ( .A(n48), .ZN(N3) );
  AOI22_X1 U76 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  INV_X1 U77 ( .A(n25), .ZN(N2) );
  AOI22_X1 U78 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_123 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n5) );
  INV_X1 U2 ( .A(n14), .ZN(n4) );
  BUF_X1 U3 ( .A(n2), .Z(n9) );
  BUF_X1 U4 ( .A(n2), .Z(n10) );
  BUF_X1 U5 ( .A(n3), .Z(n12) );
  BUF_X1 U6 ( .A(n1), .Z(n6) );
  BUF_X1 U7 ( .A(n1), .Z(n7) );
  BUF_X1 U8 ( .A(n1), .Z(n8) );
  BUF_X1 U9 ( .A(n2), .Z(n11) );
  BUF_X1 U10 ( .A(n3), .Z(n14) );
  BUF_X1 U11 ( .A(n3), .Z(n13) );
  BUF_X1 U12 ( .A(sel), .Z(n3) );
  BUF_X1 U13 ( .A(sel), .Z(n1) );
  BUF_X1 U14 ( .A(sel), .Z(n2) );
  INV_X1 U15 ( .A(n54), .ZN(N5) );
  AOI22_X1 U16 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U17 ( .A(n53), .ZN(N4) );
  AOI22_X1 U18 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U19 ( .A(n48), .ZN(N3) );
  AOI22_X1 U20 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  INV_X1 U21 ( .A(n25), .ZN(N2) );
  AOI22_X1 U22 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  INV_X1 U23 ( .A(n52), .ZN(N33) );
  AOI22_X1 U24 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n7), .ZN(n52) );
  INV_X1 U25 ( .A(n51), .ZN(N32) );
  AOI22_X1 U26 ( .A1(port0[30]), .A2(n4), .B1(port1[30]), .B2(n7), .ZN(n51) );
  INV_X1 U27 ( .A(n50), .ZN(N31) );
  AOI22_X1 U28 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  INV_X1 U29 ( .A(n49), .ZN(N30) );
  AOI22_X1 U30 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U31 ( .A(n47), .ZN(N29) );
  AOI22_X1 U32 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  INV_X1 U33 ( .A(n35), .ZN(N28) );
  AOI22_X1 U34 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  INV_X1 U35 ( .A(n33), .ZN(N27) );
  AOI22_X1 U36 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  INV_X1 U37 ( .A(n32), .ZN(N26) );
  AOI22_X1 U38 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U39 ( .A(n31), .ZN(N25) );
  AOI22_X1 U40 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  INV_X1 U41 ( .A(n30), .ZN(N24) );
  AOI22_X1 U42 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  INV_X1 U43 ( .A(n29), .ZN(N23) );
  AOI22_X1 U44 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  INV_X1 U45 ( .A(n28), .ZN(N22) );
  AOI22_X1 U46 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U47 ( .A(n27), .ZN(N21) );
  AOI22_X1 U48 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  INV_X1 U49 ( .A(n26), .ZN(N20) );
  AOI22_X1 U50 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  INV_X1 U51 ( .A(n24), .ZN(N19) );
  AOI22_X1 U52 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U53 ( .A(n23), .ZN(N18) );
  AOI22_X1 U54 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  INV_X1 U55 ( .A(n22), .ZN(N17) );
  AOI22_X1 U56 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  INV_X1 U57 ( .A(n21), .ZN(N16) );
  AOI22_X1 U58 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U59 ( .A(n20), .ZN(N15) );
  AOI22_X1 U60 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U61 ( .A(n19), .ZN(N14) );
  AOI22_X1 U62 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U63 ( .A(n18), .ZN(N13) );
  AOI22_X1 U64 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U65 ( .A(n17), .ZN(N12) );
  AOI22_X1 U66 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U67 ( .A(n16), .ZN(N11) );
  AOI22_X1 U68 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U69 ( .A(n15), .ZN(N10) );
  AOI22_X1 U70 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U71 ( .A(n58), .ZN(N9) );
  AOI22_X1 U72 ( .A1(port0[7]), .A2(n4), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U73 ( .A(n57), .ZN(N8) );
  AOI22_X1 U74 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U75 ( .A(n56), .ZN(N7) );
  AOI22_X1 U76 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U77 ( .A(n55), .ZN(N6) );
  AOI22_X1 U78 ( .A1(port0[4]), .A2(n5), .B1(port1[4]), .B2(n6), .ZN(n55) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_122 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n5) );
  INV_X1 U2 ( .A(n14), .ZN(n4) );
  BUF_X1 U3 ( .A(n2), .Z(n9) );
  BUF_X1 U4 ( .A(n2), .Z(n10) );
  BUF_X1 U5 ( .A(n3), .Z(n12) );
  BUF_X1 U6 ( .A(n1), .Z(n6) );
  BUF_X1 U7 ( .A(n1), .Z(n7) );
  BUF_X1 U8 ( .A(n1), .Z(n8) );
  BUF_X1 U9 ( .A(n2), .Z(n11) );
  BUF_X1 U10 ( .A(n3), .Z(n14) );
  BUF_X1 U11 ( .A(n3), .Z(n13) );
  BUF_X1 U12 ( .A(sel), .Z(n3) );
  BUF_X1 U13 ( .A(sel), .Z(n1) );
  BUF_X1 U14 ( .A(sel), .Z(n2) );
  INV_X1 U15 ( .A(n52), .ZN(N33) );
  AOI22_X1 U16 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n7), .ZN(n52) );
  INV_X1 U17 ( .A(n51), .ZN(N32) );
  AOI22_X1 U18 ( .A1(port0[30]), .A2(n4), .B1(port1[30]), .B2(n7), .ZN(n51) );
  INV_X1 U19 ( .A(n50), .ZN(N31) );
  AOI22_X1 U20 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  INV_X1 U21 ( .A(n49), .ZN(N30) );
  AOI22_X1 U22 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U23 ( .A(n47), .ZN(N29) );
  AOI22_X1 U24 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  INV_X1 U25 ( .A(n35), .ZN(N28) );
  AOI22_X1 U26 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  INV_X1 U27 ( .A(n33), .ZN(N27) );
  AOI22_X1 U28 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  INV_X1 U29 ( .A(n32), .ZN(N26) );
  AOI22_X1 U30 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U31 ( .A(n31), .ZN(N25) );
  AOI22_X1 U32 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  INV_X1 U33 ( .A(n30), .ZN(N24) );
  AOI22_X1 U34 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  INV_X1 U35 ( .A(n29), .ZN(N23) );
  AOI22_X1 U36 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  INV_X1 U37 ( .A(n28), .ZN(N22) );
  AOI22_X1 U38 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U39 ( .A(n27), .ZN(N21) );
  AOI22_X1 U40 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  INV_X1 U41 ( .A(n26), .ZN(N20) );
  AOI22_X1 U42 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  INV_X1 U43 ( .A(n24), .ZN(N19) );
  AOI22_X1 U44 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U45 ( .A(n23), .ZN(N18) );
  AOI22_X1 U46 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  INV_X1 U47 ( .A(n22), .ZN(N17) );
  AOI22_X1 U48 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  INV_X1 U49 ( .A(n21), .ZN(N16) );
  AOI22_X1 U50 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U51 ( .A(n20), .ZN(N15) );
  AOI22_X1 U52 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U53 ( .A(n19), .ZN(N14) );
  AOI22_X1 U54 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U55 ( .A(n18), .ZN(N13) );
  AOI22_X1 U56 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U57 ( .A(n17), .ZN(N12) );
  AOI22_X1 U58 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U59 ( .A(n16), .ZN(N11) );
  AOI22_X1 U60 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U61 ( .A(n15), .ZN(N10) );
  AOI22_X1 U62 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U63 ( .A(n57), .ZN(N8) );
  AOI22_X1 U64 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U65 ( .A(n56), .ZN(N7) );
  AOI22_X1 U66 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U67 ( .A(n55), .ZN(N6) );
  AOI22_X1 U68 ( .A1(port0[4]), .A2(n5), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U69 ( .A(n54), .ZN(N5) );
  AOI22_X1 U70 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U71 ( .A(n53), .ZN(N4) );
  AOI22_X1 U72 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U73 ( .A(n48), .ZN(N3) );
  AOI22_X1 U74 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  INV_X1 U75 ( .A(n25), .ZN(N2) );
  AOI22_X1 U76 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  INV_X1 U77 ( .A(n58), .ZN(N9) );
  AOI22_X1 U78 ( .A1(port0[7]), .A2(n5), .B1(n13), .B2(port1[7]), .ZN(n58) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_93 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  AOI22_X1 U1 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(n7), .ZN(n53) );
  AOI22_X1 U2 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  AOI22_X1 U3 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n6), .ZN(n55) );
  AOI22_X1 U4 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  AOI22_X1 U5 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n6), .ZN(n57) );
  AOI22_X1 U6 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n7), .ZN(n51) );
  AOI22_X1 U7 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n7), .ZN(n52) );
  AOI22_X1 U8 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  AOI22_X1 U9 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  AOI22_X1 U10 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  AOI22_X1 U11 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  AOI22_X1 U12 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  AOI22_X1 U13 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  AOI22_X1 U14 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  AOI22_X1 U15 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  AOI22_X1 U16 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  AOI22_X1 U17 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  AOI22_X1 U18 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  AOI22_X1 U19 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  AOI22_X1 U20 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  AOI22_X1 U21 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  AOI22_X1 U22 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  AOI22_X1 U23 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  AOI22_X1 U24 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  AOI22_X1 U25 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  AOI22_X1 U26 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  AOI22_X1 U27 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  AOI22_X1 U28 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  AOI22_X1 U29 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  AOI22_X1 U30 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  AOI22_X1 U31 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  AOI22_X1 U32 ( .A1(port0[7]), .A2(n4), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U33 ( .A(n58), .ZN(N9) );
  INV_X1 U34 ( .A(n53), .ZN(N4) );
  INV_X1 U35 ( .A(n54), .ZN(N5) );
  INV_X1 U36 ( .A(n55), .ZN(N6) );
  INV_X1 U37 ( .A(n56), .ZN(N7) );
  INV_X1 U38 ( .A(n57), .ZN(N8) );
  INV_X1 U39 ( .A(n51), .ZN(N32) );
  INV_X1 U40 ( .A(n52), .ZN(N33) );
  INV_X1 U41 ( .A(n25), .ZN(N2) );
  INV_X1 U42 ( .A(n48), .ZN(N3) );
  INV_X1 U43 ( .A(n18), .ZN(N13) );
  INV_X1 U44 ( .A(n19), .ZN(N14) );
  INV_X1 U45 ( .A(n20), .ZN(N15) );
  INV_X1 U46 ( .A(n21), .ZN(N16) );
  INV_X1 U47 ( .A(n22), .ZN(N17) );
  INV_X1 U48 ( .A(n23), .ZN(N18) );
  INV_X1 U49 ( .A(n24), .ZN(N19) );
  INV_X1 U50 ( .A(n26), .ZN(N20) );
  INV_X1 U51 ( .A(n27), .ZN(N21) );
  INV_X1 U52 ( .A(n28), .ZN(N22) );
  INV_X1 U53 ( .A(n29), .ZN(N23) );
  INV_X1 U54 ( .A(n30), .ZN(N24) );
  INV_X1 U55 ( .A(n31), .ZN(N25) );
  INV_X1 U56 ( .A(n32), .ZN(N26) );
  INV_X1 U57 ( .A(n33), .ZN(N27) );
  INV_X1 U58 ( .A(n35), .ZN(N28) );
  INV_X1 U59 ( .A(n47), .ZN(N29) );
  INV_X1 U60 ( .A(n49), .ZN(N30) );
  INV_X1 U61 ( .A(n50), .ZN(N31) );
  INV_X1 U62 ( .A(n15), .ZN(N10) );
  INV_X1 U63 ( .A(n16), .ZN(N11) );
  INV_X1 U64 ( .A(n17), .ZN(N12) );
  INV_X1 U65 ( .A(n14), .ZN(n4) );
  INV_X1 U66 ( .A(n14), .ZN(n5) );
  BUF_X1 U67 ( .A(n1), .Z(n6) );
  BUF_X1 U68 ( .A(n3), .Z(n12) );
  BUF_X1 U69 ( .A(n2), .Z(n11) );
  BUF_X1 U70 ( .A(n2), .Z(n9) );
  BUF_X1 U71 ( .A(n1), .Z(n8) );
  BUF_X1 U72 ( .A(n2), .Z(n10) );
  BUF_X1 U73 ( .A(n1), .Z(n7) );
  BUF_X1 U74 ( .A(n3), .Z(n14) );
  BUF_X1 U75 ( .A(n3), .Z(n13) );
  BUF_X1 U76 ( .A(sel), .Z(n3) );
  BUF_X1 U77 ( .A(sel), .Z(n2) );
  BUF_X1 U78 ( .A(sel), .Z(n1) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_92 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  AOI22_X1 U1 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(n7), .ZN(n53) );
  AOI22_X1 U2 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n6), .ZN(n54) );
  AOI22_X1 U3 ( .A1(port0[4]), .A2(n5), .B1(port1[4]), .B2(n6), .ZN(n55) );
  AOI22_X1 U4 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  AOI22_X1 U5 ( .A1(port0[6]), .A2(n5), .B1(port1[6]), .B2(n6), .ZN(n57) );
  AOI22_X1 U6 ( .A1(port0[30]), .A2(n4), .B1(port1[30]), .B2(n7), .ZN(n51) );
  AOI22_X1 U7 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n7), .ZN(n52) );
  AOI22_X1 U8 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  AOI22_X1 U9 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  AOI22_X1 U10 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  AOI22_X1 U11 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  AOI22_X1 U12 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  AOI22_X1 U13 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  AOI22_X1 U14 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  AOI22_X1 U15 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  AOI22_X1 U16 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  AOI22_X1 U17 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  AOI22_X1 U18 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  AOI22_X1 U19 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  AOI22_X1 U20 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  AOI22_X1 U21 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  AOI22_X1 U22 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  AOI22_X1 U23 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  AOI22_X1 U24 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  AOI22_X1 U25 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  AOI22_X1 U26 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  AOI22_X1 U27 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  AOI22_X1 U28 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  AOI22_X1 U29 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  AOI22_X1 U30 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  AOI22_X1 U31 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  AOI22_X1 U32 ( .A1(port0[7]), .A2(n4), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U33 ( .A(n58), .ZN(N9) );
  INV_X1 U34 ( .A(n53), .ZN(N4) );
  INV_X1 U35 ( .A(n54), .ZN(N5) );
  INV_X1 U36 ( .A(n55), .ZN(N6) );
  INV_X1 U37 ( .A(n56), .ZN(N7) );
  INV_X1 U38 ( .A(n57), .ZN(N8) );
  INV_X1 U39 ( .A(n51), .ZN(N32) );
  INV_X1 U40 ( .A(n52), .ZN(N33) );
  INV_X1 U41 ( .A(n25), .ZN(N2) );
  INV_X1 U42 ( .A(n48), .ZN(N3) );
  INV_X1 U43 ( .A(n18), .ZN(N13) );
  INV_X1 U44 ( .A(n19), .ZN(N14) );
  INV_X1 U45 ( .A(n20), .ZN(N15) );
  INV_X1 U46 ( .A(n21), .ZN(N16) );
  INV_X1 U47 ( .A(n22), .ZN(N17) );
  INV_X1 U48 ( .A(n23), .ZN(N18) );
  INV_X1 U49 ( .A(n24), .ZN(N19) );
  INV_X1 U50 ( .A(n26), .ZN(N20) );
  INV_X1 U51 ( .A(n27), .ZN(N21) );
  INV_X1 U52 ( .A(n28), .ZN(N22) );
  INV_X1 U53 ( .A(n29), .ZN(N23) );
  INV_X1 U54 ( .A(n30), .ZN(N24) );
  INV_X1 U55 ( .A(n31), .ZN(N25) );
  INV_X1 U56 ( .A(n32), .ZN(N26) );
  INV_X1 U57 ( .A(n33), .ZN(N27) );
  INV_X1 U58 ( .A(n35), .ZN(N28) );
  INV_X1 U59 ( .A(n47), .ZN(N29) );
  INV_X1 U60 ( .A(n49), .ZN(N30) );
  INV_X1 U61 ( .A(n50), .ZN(N31) );
  INV_X1 U62 ( .A(n15), .ZN(N10) );
  INV_X1 U63 ( .A(n16), .ZN(N11) );
  INV_X1 U64 ( .A(n17), .ZN(N12) );
  INV_X1 U65 ( .A(n14), .ZN(n4) );
  INV_X1 U66 ( .A(n14), .ZN(n5) );
  BUF_X1 U67 ( .A(n1), .Z(n6) );
  BUF_X1 U68 ( .A(n3), .Z(n12) );
  BUF_X1 U69 ( .A(n2), .Z(n11) );
  BUF_X1 U70 ( .A(n2), .Z(n9) );
  BUF_X1 U71 ( .A(n1), .Z(n8) );
  BUF_X1 U72 ( .A(n2), .Z(n10) );
  BUF_X1 U73 ( .A(n1), .Z(n7) );
  BUF_X1 U74 ( .A(n3), .Z(n14) );
  BUF_X1 U75 ( .A(n3), .Z(n13) );
  BUF_X1 U76 ( .A(sel), .Z(n3) );
  BUF_X1 U77 ( .A(sel), .Z(n2) );
  BUF_X1 U78 ( .A(sel), .Z(n1) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_91 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n58), .ZN(N9) );
  AOI22_X1 U2 ( .A1(port0[7]), .A2(n4), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U3 ( .A(n53), .ZN(N4) );
  AOI22_X1 U4 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U5 ( .A(n54), .ZN(N5) );
  AOI22_X1 U6 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U7 ( .A(n55), .ZN(N6) );
  AOI22_X1 U8 ( .A1(port0[4]), .A2(n5), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U9 ( .A(n56), .ZN(N7) );
  AOI22_X1 U10 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U11 ( .A(n57), .ZN(N8) );
  AOI22_X1 U12 ( .A1(port0[6]), .A2(n5), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U13 ( .A(n51), .ZN(N32) );
  AOI22_X1 U14 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n7), .ZN(n51) );
  INV_X1 U15 ( .A(n52), .ZN(N33) );
  AOI22_X1 U16 ( .A1(port0[31]), .A2(n4), .B1(port1[31]), .B2(n7), .ZN(n52) );
  INV_X1 U17 ( .A(n25), .ZN(N2) );
  AOI22_X1 U18 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  INV_X1 U19 ( .A(n48), .ZN(N3) );
  AOI22_X1 U20 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  INV_X1 U21 ( .A(n18), .ZN(N13) );
  AOI22_X1 U22 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U23 ( .A(n19), .ZN(N14) );
  AOI22_X1 U24 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U25 ( .A(n20), .ZN(N15) );
  AOI22_X1 U26 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U27 ( .A(n21), .ZN(N16) );
  AOI22_X1 U28 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U29 ( .A(n22), .ZN(N17) );
  AOI22_X1 U30 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  INV_X1 U31 ( .A(n23), .ZN(N18) );
  AOI22_X1 U32 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  INV_X1 U33 ( .A(n24), .ZN(N19) );
  AOI22_X1 U34 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U35 ( .A(n26), .ZN(N20) );
  AOI22_X1 U36 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  INV_X1 U37 ( .A(n27), .ZN(N21) );
  AOI22_X1 U38 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  INV_X1 U39 ( .A(n28), .ZN(N22) );
  AOI22_X1 U40 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U41 ( .A(n29), .ZN(N23) );
  AOI22_X1 U42 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  INV_X1 U43 ( .A(n30), .ZN(N24) );
  AOI22_X1 U44 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  INV_X1 U45 ( .A(n31), .ZN(N25) );
  AOI22_X1 U46 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  INV_X1 U47 ( .A(n32), .ZN(N26) );
  AOI22_X1 U48 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U49 ( .A(n33), .ZN(N27) );
  AOI22_X1 U50 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  INV_X1 U51 ( .A(n35), .ZN(N28) );
  AOI22_X1 U52 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  INV_X1 U53 ( .A(n47), .ZN(N29) );
  AOI22_X1 U54 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  INV_X1 U55 ( .A(n49), .ZN(N30) );
  AOI22_X1 U56 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U57 ( .A(n50), .ZN(N31) );
  AOI22_X1 U58 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  INV_X1 U59 ( .A(n15), .ZN(N10) );
  AOI22_X1 U60 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U61 ( .A(n16), .ZN(N11) );
  AOI22_X1 U62 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U63 ( .A(n17), .ZN(N12) );
  AOI22_X1 U64 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U65 ( .A(n14), .ZN(n4) );
  INV_X1 U66 ( .A(n14), .ZN(n5) );
  BUF_X1 U67 ( .A(n1), .Z(n6) );
  BUF_X1 U68 ( .A(n3), .Z(n12) );
  BUF_X1 U69 ( .A(n2), .Z(n11) );
  BUF_X1 U70 ( .A(n2), .Z(n9) );
  BUF_X1 U71 ( .A(n1), .Z(n8) );
  BUF_X1 U72 ( .A(n2), .Z(n10) );
  BUF_X1 U73 ( .A(n1), .Z(n7) );
  BUF_X1 U74 ( .A(n3), .Z(n14) );
  BUF_X1 U75 ( .A(n3), .Z(n13) );
  BUF_X1 U76 ( .A(sel), .Z(n3) );
  BUF_X1 U77 ( .A(sel), .Z(n2) );
  BUF_X1 U78 ( .A(sel), .Z(n1) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_90 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  BUF_X1 U3 ( .A(n1), .Z(n6) );
  BUF_X1 U4 ( .A(n3), .Z(n12) );
  BUF_X1 U5 ( .A(n2), .Z(n11) );
  BUF_X1 U6 ( .A(n2), .Z(n9) );
  BUF_X1 U7 ( .A(n1), .Z(n8) );
  BUF_X1 U8 ( .A(n2), .Z(n10) );
  BUF_X1 U9 ( .A(n1), .Z(n7) );
  BUF_X1 U10 ( .A(n3), .Z(n14) );
  BUF_X1 U11 ( .A(n3), .Z(n13) );
  BUF_X1 U12 ( .A(sel), .Z(n3) );
  BUF_X1 U13 ( .A(sel), .Z(n2) );
  BUF_X1 U14 ( .A(sel), .Z(n1) );
  INV_X1 U15 ( .A(n53), .ZN(N4) );
  AOI22_X1 U16 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U17 ( .A(n54), .ZN(N5) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U19 ( .A(n55), .ZN(N6) );
  AOI22_X1 U20 ( .A1(port0[4]), .A2(n5), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U21 ( .A(n56), .ZN(N7) );
  AOI22_X1 U22 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U23 ( .A(n57), .ZN(N8) );
  AOI22_X1 U24 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U25 ( .A(n58), .ZN(N9) );
  AOI22_X1 U26 ( .A1(port0[7]), .A2(n4), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U27 ( .A(n51), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n7), .ZN(n51) );
  INV_X1 U29 ( .A(n52), .ZN(N33) );
  AOI22_X1 U30 ( .A1(port0[31]), .A2(n4), .B1(port1[31]), .B2(n7), .ZN(n52) );
  INV_X1 U31 ( .A(n48), .ZN(N3) );
  AOI22_X1 U32 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  INV_X1 U33 ( .A(n15), .ZN(N10) );
  AOI22_X1 U34 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U35 ( .A(n16), .ZN(N11) );
  AOI22_X1 U36 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U37 ( .A(n17), .ZN(N12) );
  AOI22_X1 U38 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U39 ( .A(n18), .ZN(N13) );
  AOI22_X1 U40 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U41 ( .A(n19), .ZN(N14) );
  AOI22_X1 U42 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U43 ( .A(n20), .ZN(N15) );
  AOI22_X1 U44 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U45 ( .A(n21), .ZN(N16) );
  AOI22_X1 U46 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U47 ( .A(n22), .ZN(N17) );
  AOI22_X1 U48 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  INV_X1 U49 ( .A(n23), .ZN(N18) );
  AOI22_X1 U50 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  INV_X1 U51 ( .A(n24), .ZN(N19) );
  AOI22_X1 U52 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U53 ( .A(n26), .ZN(N20) );
  AOI22_X1 U54 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  INV_X1 U55 ( .A(n27), .ZN(N21) );
  AOI22_X1 U56 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  INV_X1 U57 ( .A(n28), .ZN(N22) );
  AOI22_X1 U58 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U59 ( .A(n29), .ZN(N23) );
  AOI22_X1 U60 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  INV_X1 U61 ( .A(n30), .ZN(N24) );
  AOI22_X1 U62 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  INV_X1 U63 ( .A(n31), .ZN(N25) );
  AOI22_X1 U64 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  INV_X1 U65 ( .A(n32), .ZN(N26) );
  AOI22_X1 U66 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U67 ( .A(n33), .ZN(N27) );
  AOI22_X1 U68 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  INV_X1 U69 ( .A(n35), .ZN(N28) );
  AOI22_X1 U70 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  INV_X1 U71 ( .A(n47), .ZN(N29) );
  AOI22_X1 U72 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  INV_X1 U73 ( .A(n49), .ZN(N30) );
  AOI22_X1 U74 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U75 ( .A(n50), .ZN(N31) );
  AOI22_X1 U76 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  INV_X1 U77 ( .A(n25), .ZN(N2) );
  AOI22_X1 U78 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_89 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  BUF_X1 U3 ( .A(n3), .Z(n14) );
  BUF_X1 U4 ( .A(n2), .Z(n11) );
  BUF_X1 U5 ( .A(n1), .Z(n8) );
  BUF_X1 U6 ( .A(n1), .Z(n7) );
  BUF_X1 U7 ( .A(n1), .Z(n6) );
  BUF_X1 U8 ( .A(n3), .Z(n13) );
  BUF_X1 U9 ( .A(n3), .Z(n12) );
  BUF_X1 U10 ( .A(n2), .Z(n10) );
  BUF_X1 U11 ( .A(n2), .Z(n9) );
  BUF_X1 U12 ( .A(sel), .Z(n3) );
  BUF_X1 U13 ( .A(sel), .Z(n2) );
  BUF_X1 U14 ( .A(sel), .Z(n1) );
  INV_X1 U15 ( .A(n25), .ZN(N2) );
  AOI22_X1 U16 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  INV_X1 U17 ( .A(n54), .ZN(N5) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U19 ( .A(n53), .ZN(N4) );
  AOI22_X1 U20 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U21 ( .A(n55), .ZN(N6) );
  AOI22_X1 U22 ( .A1(port0[4]), .A2(n5), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U23 ( .A(n56), .ZN(N7) );
  AOI22_X1 U24 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U25 ( .A(n57), .ZN(N8) );
  AOI22_X1 U26 ( .A1(port0[6]), .A2(n5), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U27 ( .A(n58), .ZN(N9) );
  AOI22_X1 U28 ( .A1(port0[7]), .A2(n5), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U29 ( .A(n48), .ZN(N3) );
  AOI22_X1 U30 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  INV_X1 U31 ( .A(n15), .ZN(N10) );
  AOI22_X1 U32 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U33 ( .A(n16), .ZN(N11) );
  AOI22_X1 U34 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U35 ( .A(n17), .ZN(N12) );
  AOI22_X1 U36 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U37 ( .A(n18), .ZN(N13) );
  AOI22_X1 U38 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U39 ( .A(n19), .ZN(N14) );
  AOI22_X1 U40 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U41 ( .A(n20), .ZN(N15) );
  AOI22_X1 U42 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U43 ( .A(n21), .ZN(N16) );
  AOI22_X1 U44 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U45 ( .A(n22), .ZN(N17) );
  AOI22_X1 U46 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  INV_X1 U47 ( .A(n23), .ZN(N18) );
  AOI22_X1 U48 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  INV_X1 U49 ( .A(n24), .ZN(N19) );
  AOI22_X1 U50 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U51 ( .A(n26), .ZN(N20) );
  AOI22_X1 U52 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  INV_X1 U53 ( .A(n27), .ZN(N21) );
  AOI22_X1 U54 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  INV_X1 U55 ( .A(n28), .ZN(N22) );
  AOI22_X1 U56 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U57 ( .A(n51), .ZN(N32) );
  AOI22_X1 U58 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n7), .ZN(n51) );
  INV_X1 U59 ( .A(n52), .ZN(N33) );
  AOI22_X1 U60 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n7), .ZN(n52) );
  INV_X1 U61 ( .A(n29), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  INV_X1 U63 ( .A(n30), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  INV_X1 U65 ( .A(n31), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  INV_X1 U67 ( .A(n32), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U69 ( .A(n33), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  INV_X1 U71 ( .A(n35), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  INV_X1 U73 ( .A(n47), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  INV_X1 U75 ( .A(n49), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U77 ( .A(n50), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_88 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X2 U1 ( .A(sel), .ZN(n1) );
  INV_X1 U2 ( .A(n28), .ZN(N4) );
  AOI22_X1 U3 ( .A1(port0[2]), .A2(n1), .B1(port1[2]), .B2(sel), .ZN(n28) );
  INV_X1 U4 ( .A(n29), .ZN(N5) );
  AOI22_X1 U5 ( .A1(port0[3]), .A2(n1), .B1(port1[3]), .B2(sel), .ZN(n29) );
  INV_X1 U6 ( .A(n30), .ZN(N6) );
  AOI22_X1 U7 ( .A1(port0[4]), .A2(n1), .B1(port1[4]), .B2(sel), .ZN(n30) );
  INV_X1 U8 ( .A(n31), .ZN(N7) );
  AOI22_X1 U9 ( .A1(port0[5]), .A2(n1), .B1(port1[5]), .B2(sel), .ZN(n31) );
  INV_X1 U10 ( .A(n32), .ZN(N8) );
  AOI22_X1 U11 ( .A1(port0[6]), .A2(n1), .B1(port1[6]), .B2(sel), .ZN(n32) );
  INV_X1 U12 ( .A(n33), .ZN(N9) );
  AOI22_X1 U13 ( .A1(port0[7]), .A2(n1), .B1(sel), .B2(port1[7]), .ZN(n33) );
  INV_X1 U14 ( .A(n26), .ZN(N32) );
  AOI22_X1 U15 ( .A1(port0[30]), .A2(n1), .B1(port1[30]), .B2(sel), .ZN(n26)
         );
  INV_X1 U16 ( .A(n27), .ZN(N33) );
  AOI22_X1 U17 ( .A1(port0[31]), .A2(n1), .B1(port1[31]), .B2(sel), .ZN(n27)
         );
  INV_X1 U18 ( .A(n23), .ZN(N3) );
  AOI22_X1 U19 ( .A1(port0[1]), .A2(n1), .B1(port1[1]), .B2(sel), .ZN(n23) );
  INV_X1 U20 ( .A(n2), .ZN(N10) );
  AOI22_X1 U21 ( .A1(port0[8]), .A2(n1), .B1(port1[8]), .B2(sel), .ZN(n2) );
  INV_X1 U22 ( .A(n3), .ZN(N11) );
  AOI22_X1 U23 ( .A1(port0[9]), .A2(n1), .B1(port1[9]), .B2(sel), .ZN(n3) );
  INV_X1 U24 ( .A(n4), .ZN(N12) );
  AOI22_X1 U25 ( .A1(port0[10]), .A2(n1), .B1(port1[10]), .B2(sel), .ZN(n4) );
  INV_X1 U26 ( .A(n5), .ZN(N13) );
  AOI22_X1 U27 ( .A1(port0[11]), .A2(n1), .B1(port1[11]), .B2(sel), .ZN(n5) );
  INV_X1 U28 ( .A(n6), .ZN(N14) );
  AOI22_X1 U29 ( .A1(port0[12]), .A2(n1), .B1(port1[12]), .B2(sel), .ZN(n6) );
  INV_X1 U30 ( .A(n7), .ZN(N15) );
  AOI22_X1 U31 ( .A1(port0[13]), .A2(n1), .B1(port1[13]), .B2(sel), .ZN(n7) );
  INV_X1 U32 ( .A(n8), .ZN(N16) );
  AOI22_X1 U33 ( .A1(port0[14]), .A2(n1), .B1(port1[14]), .B2(sel), .ZN(n8) );
  INV_X1 U34 ( .A(n9), .ZN(N17) );
  AOI22_X1 U35 ( .A1(port0[15]), .A2(n1), .B1(port1[15]), .B2(sel), .ZN(n9) );
  INV_X1 U36 ( .A(n10), .ZN(N18) );
  AOI22_X1 U37 ( .A1(port0[16]), .A2(n1), .B1(port1[16]), .B2(sel), .ZN(n10)
         );
  INV_X1 U38 ( .A(n11), .ZN(N19) );
  AOI22_X1 U39 ( .A1(port0[17]), .A2(n1), .B1(port1[17]), .B2(sel), .ZN(n11)
         );
  INV_X1 U40 ( .A(n13), .ZN(N20) );
  AOI22_X1 U41 ( .A1(port0[18]), .A2(n1), .B1(port1[18]), .B2(sel), .ZN(n13)
         );
  INV_X1 U42 ( .A(n14), .ZN(N21) );
  AOI22_X1 U43 ( .A1(port0[19]), .A2(n1), .B1(port1[19]), .B2(sel), .ZN(n14)
         );
  INV_X1 U44 ( .A(n15), .ZN(N22) );
  AOI22_X1 U45 ( .A1(port0[20]), .A2(n1), .B1(port1[20]), .B2(sel), .ZN(n15)
         );
  INV_X1 U46 ( .A(n16), .ZN(N23) );
  AOI22_X1 U47 ( .A1(port0[21]), .A2(n1), .B1(port1[21]), .B2(sel), .ZN(n16)
         );
  INV_X1 U48 ( .A(n17), .ZN(N24) );
  AOI22_X1 U49 ( .A1(port0[22]), .A2(n1), .B1(port1[22]), .B2(sel), .ZN(n17)
         );
  INV_X1 U50 ( .A(n18), .ZN(N25) );
  AOI22_X1 U51 ( .A1(port0[23]), .A2(n1), .B1(port1[23]), .B2(sel), .ZN(n18)
         );
  INV_X1 U52 ( .A(n19), .ZN(N26) );
  AOI22_X1 U53 ( .A1(port0[24]), .A2(n1), .B1(port1[24]), .B2(sel), .ZN(n19)
         );
  INV_X1 U54 ( .A(n20), .ZN(N27) );
  AOI22_X1 U55 ( .A1(port0[25]), .A2(n1), .B1(port1[25]), .B2(sel), .ZN(n20)
         );
  INV_X1 U56 ( .A(n21), .ZN(N28) );
  AOI22_X1 U57 ( .A1(port0[26]), .A2(n1), .B1(port1[26]), .B2(sel), .ZN(n21)
         );
  INV_X1 U58 ( .A(n22), .ZN(N29) );
  AOI22_X1 U59 ( .A1(port0[27]), .A2(n1), .B1(port1[27]), .B2(sel), .ZN(n22)
         );
  INV_X1 U60 ( .A(n24), .ZN(N30) );
  AOI22_X1 U61 ( .A1(port0[28]), .A2(n1), .B1(port1[28]), .B2(sel), .ZN(n24)
         );
  INV_X1 U62 ( .A(n25), .ZN(N31) );
  AOI22_X1 U63 ( .A1(port0[29]), .A2(n1), .B1(port1[29]), .B2(sel), .ZN(n25)
         );
  INV_X1 U64 ( .A(n12), .ZN(N2) );
  AOI22_X1 U65 ( .A1(port0[0]), .A2(n1), .B1(port1[0]), .B2(sel), .ZN(n12) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_87 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n37, n38;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n4), .ZN(n1) );
  INV_X1 U2 ( .A(n4), .ZN(n2) );
  BUF_X1 U3 ( .A(sel), .Z(n4) );
  BUF_X1 U4 ( .A(sel), .Z(n3) );
  INV_X1 U5 ( .A(n29), .ZN(N32) );
  AOI22_X1 U6 ( .A1(port0[30]), .A2(n2), .B1(port1[30]), .B2(sel), .ZN(n29) );
  INV_X1 U7 ( .A(n28), .ZN(N31) );
  AOI22_X1 U8 ( .A1(port0[29]), .A2(n2), .B1(port1[29]), .B2(sel), .ZN(n28) );
  INV_X1 U9 ( .A(n27), .ZN(N30) );
  AOI22_X1 U10 ( .A1(port0[28]), .A2(n2), .B1(port1[28]), .B2(sel), .ZN(n27)
         );
  INV_X1 U11 ( .A(n25), .ZN(N29) );
  AOI22_X1 U12 ( .A1(port0[27]), .A2(n2), .B1(port1[27]), .B2(sel), .ZN(n25)
         );
  INV_X1 U13 ( .A(n24), .ZN(N28) );
  AOI22_X1 U14 ( .A1(port0[26]), .A2(n2), .B1(port1[26]), .B2(sel), .ZN(n24)
         );
  AOI22_X1 U15 ( .A1(port0[31]), .A2(n2), .B1(port1[31]), .B2(sel), .ZN(n30)
         );
  INV_X1 U16 ( .A(n31), .ZN(N4) );
  AOI22_X1 U17 ( .A1(port0[2]), .A2(n1), .B1(port1[2]), .B2(sel), .ZN(n31) );
  INV_X1 U18 ( .A(n32), .ZN(N5) );
  AOI22_X1 U19 ( .A1(port0[3]), .A2(n2), .B1(port1[3]), .B2(sel), .ZN(n32) );
  INV_X1 U20 ( .A(n33), .ZN(N6) );
  AOI22_X1 U21 ( .A1(port0[4]), .A2(n1), .B1(port1[4]), .B2(sel), .ZN(n33) );
  INV_X1 U22 ( .A(n35), .ZN(N7) );
  AOI22_X1 U23 ( .A1(port0[5]), .A2(n2), .B1(port1[5]), .B2(sel), .ZN(n35) );
  INV_X1 U24 ( .A(n37), .ZN(N8) );
  AOI22_X1 U25 ( .A1(port0[6]), .A2(n1), .B1(port1[6]), .B2(sel), .ZN(n37) );
  INV_X1 U26 ( .A(n38), .ZN(N9) );
  AOI22_X1 U27 ( .A1(port0[7]), .A2(n1), .B1(n3), .B2(port1[7]), .ZN(n38) );
  INV_X1 U28 ( .A(n23), .ZN(N27) );
  AOI22_X1 U29 ( .A1(port0[25]), .A2(n2), .B1(port1[25]), .B2(sel), .ZN(n23)
         );
  INV_X1 U30 ( .A(n22), .ZN(N26) );
  AOI22_X1 U31 ( .A1(port0[24]), .A2(n2), .B1(port1[24]), .B2(sel), .ZN(n22)
         );
  INV_X1 U32 ( .A(n21), .ZN(N25) );
  AOI22_X1 U33 ( .A1(port0[23]), .A2(n2), .B1(port1[23]), .B2(sel), .ZN(n21)
         );
  INV_X1 U34 ( .A(n20), .ZN(N24) );
  AOI22_X1 U35 ( .A1(port0[22]), .A2(n2), .B1(port1[22]), .B2(sel), .ZN(n20)
         );
  INV_X1 U36 ( .A(n19), .ZN(N23) );
  AOI22_X1 U37 ( .A1(port0[21]), .A2(n2), .B1(port1[21]), .B2(sel), .ZN(n19)
         );
  INV_X1 U38 ( .A(n18), .ZN(N22) );
  AOI22_X1 U39 ( .A1(port0[20]), .A2(n2), .B1(port1[20]), .B2(sel), .ZN(n18)
         );
  INV_X1 U40 ( .A(n17), .ZN(N21) );
  AOI22_X1 U41 ( .A1(port0[19]), .A2(n2), .B1(port1[19]), .B2(sel), .ZN(n17)
         );
  INV_X1 U42 ( .A(n16), .ZN(N20) );
  AOI22_X1 U43 ( .A1(port0[18]), .A2(n1), .B1(port1[18]), .B2(sel), .ZN(n16)
         );
  INV_X1 U44 ( .A(n9), .ZN(N14) );
  AOI22_X1 U45 ( .A1(port0[12]), .A2(n1), .B1(port1[12]), .B2(sel), .ZN(n9) );
  INV_X1 U46 ( .A(n10), .ZN(N15) );
  AOI22_X1 U47 ( .A1(port0[13]), .A2(n1), .B1(port1[13]), .B2(n3), .ZN(n10) );
  INV_X1 U48 ( .A(n11), .ZN(N16) );
  AOI22_X1 U49 ( .A1(port0[14]), .A2(n1), .B1(port1[14]), .B2(n3), .ZN(n11) );
  INV_X1 U50 ( .A(n14), .ZN(N19) );
  AOI22_X1 U51 ( .A1(port0[17]), .A2(n1), .B1(port1[17]), .B2(sel), .ZN(n14)
         );
  INV_X1 U52 ( .A(n13), .ZN(N18) );
  AOI22_X1 U53 ( .A1(port0[16]), .A2(n1), .B1(port1[16]), .B2(sel), .ZN(n13)
         );
  INV_X1 U54 ( .A(n12), .ZN(N17) );
  AOI22_X1 U55 ( .A1(port0[15]), .A2(n1), .B1(port1[15]), .B2(sel), .ZN(n12)
         );
  INV_X1 U56 ( .A(n15), .ZN(N2) );
  AOI22_X1 U57 ( .A1(port0[0]), .A2(n1), .B1(port1[0]), .B2(sel), .ZN(n15) );
  INV_X1 U58 ( .A(n26), .ZN(N3) );
  AOI22_X1 U59 ( .A1(port0[1]), .A2(n2), .B1(port1[1]), .B2(sel), .ZN(n26) );
  INV_X1 U60 ( .A(n5), .ZN(N10) );
  AOI22_X1 U61 ( .A1(port0[8]), .A2(n1), .B1(port1[8]), .B2(n3), .ZN(n5) );
  INV_X1 U62 ( .A(n6), .ZN(N11) );
  AOI22_X1 U63 ( .A1(port0[9]), .A2(n1), .B1(port1[9]), .B2(n3), .ZN(n6) );
  INV_X1 U64 ( .A(n7), .ZN(N12) );
  AOI22_X1 U65 ( .A1(port0[10]), .A2(n1), .B1(port1[10]), .B2(n3), .ZN(n7) );
  INV_X1 U66 ( .A(n8), .ZN(N13) );
  AOI22_X1 U67 ( .A1(port0[11]), .A2(n1), .B1(port1[11]), .B2(sel), .ZN(n8) );
  INV_X1 U68 ( .A(n30), .ZN(N33) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_86 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n39, n40, n41, n42;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n6), .ZN(n1) );
  INV_X1 U2 ( .A(n6), .ZN(n2) );
  BUF_X1 U3 ( .A(sel), .Z(n3) );
  BUF_X1 U4 ( .A(sel), .Z(n4) );
  BUF_X1 U5 ( .A(n4), .Z(n6) );
  BUF_X1 U6 ( .A(n3), .Z(n5) );
  INV_X1 U7 ( .A(n31), .ZN(N32) );
  AOI22_X1 U8 ( .A1(port0[30]), .A2(n2), .B1(port1[30]), .B2(n4), .ZN(n31) );
  INV_X1 U9 ( .A(n30), .ZN(N31) );
  AOI22_X1 U10 ( .A1(port0[29]), .A2(n2), .B1(port1[29]), .B2(n3), .ZN(n30) );
  INV_X1 U11 ( .A(n29), .ZN(N30) );
  AOI22_X1 U12 ( .A1(port0[28]), .A2(n2), .B1(port1[28]), .B2(n4), .ZN(n29) );
  INV_X1 U13 ( .A(n27), .ZN(N29) );
  AOI22_X1 U14 ( .A1(port0[27]), .A2(n2), .B1(port1[27]), .B2(n4), .ZN(n27) );
  INV_X1 U15 ( .A(n26), .ZN(N28) );
  AOI22_X1 U16 ( .A1(port0[26]), .A2(n2), .B1(port1[26]), .B2(n4), .ZN(n26) );
  INV_X1 U17 ( .A(n32), .ZN(N33) );
  INV_X1 U18 ( .A(n33), .ZN(N4) );
  AOI22_X1 U19 ( .A1(port0[2]), .A2(n2), .B1(port1[2]), .B2(n4), .ZN(n33) );
  INV_X1 U20 ( .A(n35), .ZN(N5) );
  AOI22_X1 U21 ( .A1(port0[3]), .A2(n1), .B1(port1[3]), .B2(n3), .ZN(n35) );
  INV_X1 U22 ( .A(n39), .ZN(N6) );
  AOI22_X1 U23 ( .A1(port0[4]), .A2(n2), .B1(port1[4]), .B2(n3), .ZN(n39) );
  INV_X1 U24 ( .A(n40), .ZN(N7) );
  AOI22_X1 U25 ( .A1(port0[5]), .A2(n1), .B1(port1[5]), .B2(n3), .ZN(n40) );
  INV_X1 U26 ( .A(n41), .ZN(N8) );
  AOI22_X1 U27 ( .A1(port0[6]), .A2(n2), .B1(port1[6]), .B2(n3), .ZN(n41) );
  INV_X1 U28 ( .A(n42), .ZN(N9) );
  AOI22_X1 U29 ( .A1(port0[7]), .A2(n1), .B1(n5), .B2(port1[7]), .ZN(n42) );
  INV_X1 U30 ( .A(n25), .ZN(N27) );
  AOI22_X1 U31 ( .A1(port0[25]), .A2(n2), .B1(port1[25]), .B2(n4), .ZN(n25) );
  INV_X1 U32 ( .A(n24), .ZN(N26) );
  AOI22_X1 U33 ( .A1(port0[24]), .A2(n2), .B1(port1[24]), .B2(n4), .ZN(n24) );
  INV_X1 U34 ( .A(n23), .ZN(N25) );
  AOI22_X1 U35 ( .A1(port0[23]), .A2(n2), .B1(port1[23]), .B2(n3), .ZN(n23) );
  INV_X1 U36 ( .A(n22), .ZN(N24) );
  AOI22_X1 U37 ( .A1(port0[22]), .A2(n2), .B1(port1[22]), .B2(n4), .ZN(n22) );
  INV_X1 U38 ( .A(n21), .ZN(N23) );
  AOI22_X1 U39 ( .A1(port0[21]), .A2(n2), .B1(port1[21]), .B2(n3), .ZN(n21) );
  INV_X1 U40 ( .A(n20), .ZN(N22) );
  AOI22_X1 U41 ( .A1(port0[20]), .A2(n2), .B1(port1[20]), .B2(n4), .ZN(n20) );
  INV_X1 U42 ( .A(n19), .ZN(N21) );
  AOI22_X1 U43 ( .A1(port0[19]), .A2(n2), .B1(port1[19]), .B2(n3), .ZN(n19) );
  INV_X1 U44 ( .A(n18), .ZN(N20) );
  AOI22_X1 U45 ( .A1(port0[18]), .A2(n1), .B1(port1[18]), .B2(n4), .ZN(n18) );
  INV_X1 U46 ( .A(n11), .ZN(N14) );
  AOI22_X1 U47 ( .A1(port0[12]), .A2(n1), .B1(port1[12]), .B2(n3), .ZN(n11) );
  INV_X1 U48 ( .A(n12), .ZN(N15) );
  AOI22_X1 U49 ( .A1(port0[13]), .A2(n1), .B1(port1[13]), .B2(n5), .ZN(n12) );
  INV_X1 U50 ( .A(n13), .ZN(N16) );
  AOI22_X1 U51 ( .A1(port0[14]), .A2(n1), .B1(port1[14]), .B2(n5), .ZN(n13) );
  INV_X1 U52 ( .A(n16), .ZN(N19) );
  AOI22_X1 U53 ( .A1(port0[17]), .A2(n1), .B1(port1[17]), .B2(n4), .ZN(n16) );
  INV_X1 U54 ( .A(n15), .ZN(N18) );
  AOI22_X1 U55 ( .A1(port0[16]), .A2(n1), .B1(port1[16]), .B2(n3), .ZN(n15) );
  INV_X1 U56 ( .A(n14), .ZN(N17) );
  AOI22_X1 U57 ( .A1(port0[15]), .A2(n1), .B1(port1[15]), .B2(n3), .ZN(n14) );
  INV_X1 U58 ( .A(n17), .ZN(N2) );
  AOI22_X1 U59 ( .A1(port0[0]), .A2(n1), .B1(port1[0]), .B2(n4), .ZN(n17) );
  INV_X1 U60 ( .A(n28), .ZN(N3) );
  AOI22_X1 U61 ( .A1(port0[1]), .A2(n2), .B1(port1[1]), .B2(n4), .ZN(n28) );
  INV_X1 U62 ( .A(n7), .ZN(N10) );
  AOI22_X1 U63 ( .A1(port0[8]), .A2(n1), .B1(port1[8]), .B2(n5), .ZN(n7) );
  INV_X1 U64 ( .A(n8), .ZN(N11) );
  AOI22_X1 U65 ( .A1(port0[9]), .A2(n1), .B1(port1[9]), .B2(n5), .ZN(n8) );
  INV_X1 U66 ( .A(n9), .ZN(N12) );
  AOI22_X1 U67 ( .A1(port0[10]), .A2(n1), .B1(port1[10]), .B2(n5), .ZN(n9) );
  INV_X1 U68 ( .A(n10), .ZN(N13) );
  AOI22_X1 U69 ( .A1(port0[11]), .A2(n1), .B1(port1[11]), .B2(n4), .ZN(n10) );
  AOI22_X1 U70 ( .A1(port0[31]), .A2(n1), .B1(port1[31]), .B2(n4), .ZN(n32) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_85 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n5) );
  INV_X1 U2 ( .A(n14), .ZN(n4) );
  BUF_X1 U3 ( .A(n1), .Z(n6) );
  BUF_X1 U4 ( .A(n1), .Z(n7) );
  BUF_X1 U5 ( .A(n2), .Z(n9) );
  BUF_X1 U6 ( .A(n2), .Z(n10) );
  BUF_X1 U7 ( .A(n1), .Z(n8) );
  BUF_X1 U8 ( .A(n3), .Z(n12) );
  BUF_X1 U9 ( .A(n2), .Z(n11) );
  BUF_X1 U10 ( .A(n3), .Z(n14) );
  BUF_X1 U11 ( .A(n3), .Z(n13) );
  AOI22_X1 U12 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n6), .ZN(n57) );
  AOI22_X1 U13 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  AOI22_X1 U14 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n6), .ZN(n55) );
  AOI22_X1 U15 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  AOI22_X1 U16 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n7), .ZN(n53) );
  AOI22_X1 U17 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n7), .ZN(n51) );
  AOI22_X1 U18 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  AOI22_X1 U19 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  AOI22_X1 U20 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  AOI22_X1 U21 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  AOI22_X1 U22 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  AOI22_X1 U23 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  AOI22_X1 U24 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  AOI22_X1 U25 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  AOI22_X1 U26 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  AOI22_X1 U27 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  AOI22_X1 U28 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  AOI22_X1 U29 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  AOI22_X1 U30 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  AOI22_X1 U31 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  AOI22_X1 U32 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  INV_X1 U33 ( .A(n58), .ZN(N9) );
  AOI22_X1 U34 ( .A1(port0[7]), .A2(n5), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U35 ( .A(n32), .ZN(N26) );
  AOI22_X1 U36 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U37 ( .A(n17), .ZN(N12) );
  AOI22_X1 U38 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U39 ( .A(n19), .ZN(N14) );
  AOI22_X1 U40 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U41 ( .A(n49), .ZN(N30) );
  AOI22_X1 U42 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U43 ( .A(n28), .ZN(N22) );
  AOI22_X1 U44 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U45 ( .A(n24), .ZN(N19) );
  AOI22_X1 U46 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U47 ( .A(n20), .ZN(N15) );
  AOI22_X1 U48 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U49 ( .A(n18), .ZN(N13) );
  AOI22_X1 U50 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U51 ( .A(n25), .ZN(N2) );
  AOI22_X1 U52 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  INV_X1 U53 ( .A(n52), .ZN(N33) );
  AOI22_X1 U54 ( .A1(port0[31]), .A2(n4), .B1(port1[31]), .B2(n7), .ZN(n52) );
  BUF_X1 U55 ( .A(sel), .Z(n3) );
  BUF_X1 U56 ( .A(sel), .Z(n1) );
  BUF_X1 U57 ( .A(sel), .Z(n2) );
  INV_X1 U58 ( .A(n57), .ZN(N8) );
  INV_X1 U59 ( .A(n54), .ZN(N5) );
  INV_X1 U60 ( .A(n55), .ZN(N6) );
  INV_X1 U61 ( .A(n56), .ZN(N7) );
  INV_X1 U62 ( .A(n53), .ZN(N4) );
  INV_X1 U63 ( .A(n51), .ZN(N32) );
  INV_X1 U64 ( .A(n15), .ZN(N10) );
  INV_X1 U65 ( .A(n16), .ZN(N11) );
  INV_X1 U66 ( .A(n50), .ZN(N31) );
  INV_X1 U67 ( .A(n35), .ZN(N28) );
  INV_X1 U68 ( .A(n29), .ZN(N23) );
  INV_X1 U69 ( .A(n30), .ZN(N24) );
  INV_X1 U70 ( .A(n31), .ZN(N25) );
  INV_X1 U71 ( .A(n26), .ZN(N20) );
  INV_X1 U72 ( .A(n27), .ZN(N21) );
  INV_X1 U73 ( .A(n48), .ZN(N3) );
  INV_X1 U74 ( .A(n21), .ZN(N16) );
  INV_X1 U75 ( .A(n22), .ZN(N17) );
  INV_X1 U76 ( .A(n23), .ZN(N18) );
  INV_X1 U77 ( .A(n33), .ZN(N27) );
  INV_X1 U78 ( .A(n47), .ZN(N29) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_84 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n5) );
  INV_X1 U2 ( .A(n14), .ZN(n4) );
  BUF_X1 U3 ( .A(n1), .Z(n6) );
  BUF_X1 U4 ( .A(n2), .Z(n9) );
  BUF_X1 U5 ( .A(n2), .Z(n10) );
  BUF_X1 U6 ( .A(n1), .Z(n8) );
  BUF_X1 U7 ( .A(n3), .Z(n12) );
  BUF_X1 U8 ( .A(n2), .Z(n11) );
  BUF_X1 U9 ( .A(n3), .Z(n14) );
  BUF_X1 U10 ( .A(n3), .Z(n13) );
  BUF_X1 U11 ( .A(n1), .Z(n7) );
  BUF_X1 U12 ( .A(sel), .Z(n3) );
  BUF_X1 U13 ( .A(sel), .Z(n1) );
  BUF_X1 U14 ( .A(sel), .Z(n2) );
  INV_X1 U15 ( .A(n57), .ZN(N8) );
  AOI22_X1 U16 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U17 ( .A(n54), .ZN(N5) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U19 ( .A(n55), .ZN(N6) );
  AOI22_X1 U20 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U21 ( .A(n56), .ZN(N7) );
  AOI22_X1 U22 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U23 ( .A(n53), .ZN(N4) );
  AOI22_X1 U24 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U25 ( .A(n51), .ZN(N32) );
  AOI22_X1 U26 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n7), .ZN(n51) );
  INV_X1 U27 ( .A(n15), .ZN(N10) );
  AOI22_X1 U28 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U29 ( .A(n16), .ZN(N11) );
  AOI22_X1 U30 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U31 ( .A(n50), .ZN(N31) );
  AOI22_X1 U32 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  INV_X1 U33 ( .A(n35), .ZN(N28) );
  AOI22_X1 U34 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  INV_X1 U35 ( .A(n29), .ZN(N23) );
  AOI22_X1 U36 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  INV_X1 U37 ( .A(n30), .ZN(N24) );
  AOI22_X1 U38 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  INV_X1 U39 ( .A(n31), .ZN(N25) );
  AOI22_X1 U40 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  INV_X1 U41 ( .A(n26), .ZN(N20) );
  AOI22_X1 U42 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  INV_X1 U43 ( .A(n27), .ZN(N21) );
  AOI22_X1 U44 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  INV_X1 U45 ( .A(n48), .ZN(N3) );
  AOI22_X1 U46 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  INV_X1 U47 ( .A(n21), .ZN(N16) );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U49 ( .A(n22), .ZN(N17) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  INV_X1 U51 ( .A(n23), .ZN(N18) );
  AOI22_X1 U52 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  INV_X1 U53 ( .A(n28), .ZN(N22) );
  AOI22_X1 U54 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U55 ( .A(n24), .ZN(N19) );
  AOI22_X1 U56 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U57 ( .A(n20), .ZN(N15) );
  AOI22_X1 U58 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U59 ( .A(n25), .ZN(N2) );
  AOI22_X1 U60 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  INV_X1 U61 ( .A(n52), .ZN(N33) );
  INV_X1 U62 ( .A(n49), .ZN(N30) );
  AOI22_X1 U63 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U64 ( .A(n32), .ZN(N26) );
  AOI22_X1 U65 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U66 ( .A(n58), .ZN(N9) );
  AOI22_X1 U67 ( .A1(port0[7]), .A2(n5), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U68 ( .A(n17), .ZN(N12) );
  AOI22_X1 U69 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U70 ( .A(n18), .ZN(N13) );
  AOI22_X1 U71 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U72 ( .A(n19), .ZN(N14) );
  AOI22_X1 U73 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U74 ( .A(n33), .ZN(N27) );
  AOI22_X1 U75 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  INV_X1 U76 ( .A(n47), .ZN(N29) );
  AOI22_X1 U77 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  AOI22_X1 U78 ( .A1(port0[31]), .A2(n4), .B1(port1[31]), .B2(n7), .ZN(n52) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_83 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  CLKBUF_X1 U1 ( .A(n3), .Z(n14) );
  BUF_X1 U2 ( .A(n2), .Z(n10) );
  BUF_X1 U3 ( .A(n3), .Z(n15) );
  INV_X1 U4 ( .A(n15), .ZN(n4) );
  INV_X1 U5 ( .A(n15), .ZN(n5) );
  INV_X1 U6 ( .A(n57), .ZN(N6) );
  INV_X1 U7 ( .A(n53), .ZN(N32) );
  INV_X1 U8 ( .A(n59), .ZN(N8) );
  INV_X1 U9 ( .A(n58), .ZN(N7) );
  INV_X1 U10 ( .A(n26), .ZN(N2) );
  INV_X1 U11 ( .A(n17), .ZN(N11) );
  INV_X1 U12 ( .A(n35), .ZN(N27) );
  INV_X1 U13 ( .A(n51), .ZN(N30) );
  INV_X1 U14 ( .A(n29), .ZN(N22) );
  INV_X1 U15 ( .A(n48), .ZN(N28) );
  INV_X1 U16 ( .A(n50), .ZN(N3) );
  INV_X1 U17 ( .A(n52), .ZN(N31) );
  INV_X1 U18 ( .A(n49), .ZN(N29) );
  INV_X1 U19 ( .A(n23), .ZN(N17) );
  INV_X1 U20 ( .A(n18), .ZN(N12) );
  INV_X1 U21 ( .A(n20), .ZN(N14) );
  INV_X1 U22 ( .A(n30), .ZN(N23) );
  INV_X1 U23 ( .A(n16), .ZN(N10) );
  INV_X1 U24 ( .A(n32), .ZN(N25) );
  INV_X1 U25 ( .A(n19), .ZN(N13) );
  INV_X1 U26 ( .A(n27), .ZN(N20) );
  INV_X1 U27 ( .A(n31), .ZN(N24) );
  INV_X1 U28 ( .A(n24), .ZN(N18) );
  INV_X1 U29 ( .A(n21), .ZN(N15) );
  INV_X1 U30 ( .A(n60), .ZN(N9) );
  INV_X1 U31 ( .A(n54), .ZN(N33) );
  INV_X1 U32 ( .A(n55), .ZN(N4) );
  INV_X1 U33 ( .A(n56), .ZN(N5) );
  BUF_X1 U34 ( .A(n1), .Z(n8) );
  CLKBUF_X1 U35 ( .A(n1), .Z(n7) );
  BUF_X1 U36 ( .A(n2), .Z(n12) );
  CLKBUF_X1 U37 ( .A(n2), .Z(n11) );
  CLKBUF_X1 U38 ( .A(n1), .Z(n9) );
  BUF_X1 U39 ( .A(n3), .Z(n13) );
  INV_X1 U40 ( .A(n22), .ZN(N16) );
  INV_X1 U41 ( .A(n25), .ZN(N19) );
  INV_X1 U42 ( .A(n28), .ZN(N21) );
  INV_X1 U43 ( .A(n33), .ZN(N26) );
  AOI22_X1 U44 ( .A1(port0[4]), .A2(n6), .B1(port1[4]), .B2(n7), .ZN(n57) );
  AOI22_X1 U45 ( .A1(port0[31]), .A2(n6), .B1(port1[31]), .B2(n8), .ZN(n54) );
  AOI22_X1 U46 ( .A1(port0[2]), .A2(n6), .B1(port1[2]), .B2(n8), .ZN(n55) );
  AOI22_X1 U47 ( .A1(port0[3]), .A2(n6), .B1(port1[3]), .B2(n7), .ZN(n56) );
  AOI22_X1 U48 ( .A1(port0[30]), .A2(n6), .B1(port1[30]), .B2(n8), .ZN(n53) );
  AOI22_X1 U49 ( .A1(port0[7]), .A2(n6), .B1(n14), .B2(port1[7]), .ZN(n60) );
  AOI22_X1 U50 ( .A1(port0[6]), .A2(n6), .B1(port1[6]), .B2(n7), .ZN(n59) );
  AOI22_X1 U51 ( .A1(port0[5]), .A2(n6), .B1(port1[5]), .B2(n7), .ZN(n58) );
  AOI22_X1 U52 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n12), .ZN(n26) );
  AOI22_X1 U53 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n9), .ZN(n48) );
  AOI22_X1 U54 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U55 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n9), .ZN(n50) );
  AOI22_X1 U56 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n9), .ZN(n35) );
  AOI22_X1 U57 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n14), .ZN(n17) );
  AOI22_X1 U58 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n10), .ZN(n32)
         );
  AOI22_X1 U59 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n14), .ZN(n16) );
  AOI22_X1 U60 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n13), .ZN(n22)
         );
  AOI22_X1 U61 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n9), .ZN(n49) );
  AOI22_X1 U62 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n10), .ZN(n31)
         );
  AOI22_X1 U63 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n14), .ZN(n18)
         );
  AOI22_X1 U64 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n13), .ZN(n19)
         );
  AOI22_X1 U65 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n8), .ZN(n51) );
  AOI22_X1 U66 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n12), .ZN(n23)
         );
  AOI22_X1 U67 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n11), .ZN(n28)
         );
  AOI22_X1 U68 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n11), .ZN(n27)
         );
  AOI22_X1 U69 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n10), .ZN(n30)
         );
  AOI22_X1 U70 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n13), .ZN(n20)
         );
  AOI22_X1 U71 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n12), .ZN(n25)
         );
  AOI22_X1 U72 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n13), .ZN(n21)
         );
  AOI22_X1 U73 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n12), .ZN(n24)
         );
  AOI22_X1 U74 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n10), .ZN(n33)
         );
  AOI22_X1 U75 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n11), .ZN(n29)
         );
  CLKBUF_X1 U76 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U77 ( .A(sel), .Z(n1) );
  CLKBUF_X1 U78 ( .A(sel), .Z(n2) );
  INV_X1 U79 ( .A(n15), .ZN(n6) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_82 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  CLKBUF_X1 U1 ( .A(n3), .Z(n14) );
  BUF_X1 U2 ( .A(n2), .Z(n10) );
  BUF_X1 U3 ( .A(n3), .Z(n15) );
  INV_X1 U4 ( .A(n15), .ZN(n4) );
  INV_X1 U5 ( .A(n15), .ZN(n5) );
  INV_X1 U6 ( .A(n57), .ZN(N6) );
  INV_X1 U7 ( .A(n53), .ZN(N32) );
  INV_X1 U8 ( .A(n59), .ZN(N8) );
  INV_X1 U9 ( .A(n58), .ZN(N7) );
  INV_X1 U10 ( .A(n26), .ZN(N2) );
  INV_X1 U11 ( .A(n17), .ZN(N11) );
  INV_X1 U12 ( .A(n35), .ZN(N27) );
  INV_X1 U13 ( .A(n51), .ZN(N30) );
  INV_X1 U14 ( .A(n29), .ZN(N22) );
  INV_X1 U15 ( .A(n48), .ZN(N28) );
  INV_X1 U16 ( .A(n50), .ZN(N3) );
  INV_X1 U17 ( .A(n52), .ZN(N31) );
  INV_X1 U18 ( .A(n49), .ZN(N29) );
  INV_X1 U19 ( .A(n23), .ZN(N17) );
  INV_X1 U20 ( .A(n18), .ZN(N12) );
  INV_X1 U21 ( .A(n20), .ZN(N14) );
  INV_X1 U22 ( .A(n30), .ZN(N23) );
  INV_X1 U23 ( .A(n16), .ZN(N10) );
  INV_X1 U24 ( .A(n32), .ZN(N25) );
  INV_X1 U25 ( .A(n19), .ZN(N13) );
  INV_X1 U26 ( .A(n27), .ZN(N20) );
  INV_X1 U27 ( .A(n31), .ZN(N24) );
  INV_X1 U28 ( .A(n24), .ZN(N18) );
  INV_X1 U29 ( .A(n21), .ZN(N15) );
  INV_X1 U30 ( .A(n60), .ZN(N9) );
  INV_X1 U31 ( .A(n54), .ZN(N33) );
  INV_X1 U32 ( .A(n55), .ZN(N4) );
  INV_X1 U33 ( .A(n56), .ZN(N5) );
  BUF_X1 U34 ( .A(n1), .Z(n8) );
  CLKBUF_X1 U35 ( .A(n1), .Z(n7) );
  BUF_X1 U36 ( .A(n2), .Z(n12) );
  CLKBUF_X1 U37 ( .A(n2), .Z(n11) );
  CLKBUF_X1 U38 ( .A(n1), .Z(n9) );
  BUF_X1 U39 ( .A(n3), .Z(n13) );
  INV_X1 U40 ( .A(n22), .ZN(N16) );
  INV_X1 U41 ( .A(n25), .ZN(N19) );
  INV_X1 U42 ( .A(n28), .ZN(N21) );
  INV_X1 U43 ( .A(n33), .ZN(N26) );
  AOI22_X1 U44 ( .A1(port0[4]), .A2(n6), .B1(port1[4]), .B2(n7), .ZN(n57) );
  AOI22_X1 U45 ( .A1(port0[31]), .A2(n6), .B1(port1[31]), .B2(n8), .ZN(n54) );
  AOI22_X1 U46 ( .A1(port0[2]), .A2(n6), .B1(port1[2]), .B2(n8), .ZN(n55) );
  AOI22_X1 U47 ( .A1(port0[3]), .A2(n6), .B1(port1[3]), .B2(n7), .ZN(n56) );
  AOI22_X1 U48 ( .A1(port0[30]), .A2(n6), .B1(port1[30]), .B2(n8), .ZN(n53) );
  AOI22_X1 U49 ( .A1(port0[7]), .A2(n6), .B1(n14), .B2(port1[7]), .ZN(n60) );
  AOI22_X1 U50 ( .A1(port0[6]), .A2(n6), .B1(port1[6]), .B2(n7), .ZN(n59) );
  AOI22_X1 U51 ( .A1(port0[5]), .A2(n6), .B1(port1[5]), .B2(n7), .ZN(n58) );
  AOI22_X1 U52 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n12), .ZN(n26) );
  AOI22_X1 U53 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n9), .ZN(n48) );
  AOI22_X1 U54 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U55 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n9), .ZN(n50) );
  AOI22_X1 U56 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n9), .ZN(n35) );
  AOI22_X1 U57 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n14), .ZN(n17) );
  AOI22_X1 U58 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n10), .ZN(n32)
         );
  AOI22_X1 U59 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n14), .ZN(n16) );
  AOI22_X1 U60 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n13), .ZN(n22)
         );
  AOI22_X1 U61 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n9), .ZN(n49) );
  AOI22_X1 U62 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n10), .ZN(n31)
         );
  AOI22_X1 U63 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n14), .ZN(n18)
         );
  AOI22_X1 U64 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n13), .ZN(n19)
         );
  AOI22_X1 U65 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n8), .ZN(n51) );
  AOI22_X1 U66 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n12), .ZN(n23)
         );
  AOI22_X1 U67 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n11), .ZN(n28)
         );
  AOI22_X1 U68 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n11), .ZN(n27)
         );
  AOI22_X1 U69 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n10), .ZN(n30)
         );
  AOI22_X1 U70 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n13), .ZN(n20)
         );
  AOI22_X1 U71 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n12), .ZN(n25)
         );
  AOI22_X1 U72 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n13), .ZN(n21)
         );
  AOI22_X1 U73 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n12), .ZN(n24)
         );
  AOI22_X1 U74 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n10), .ZN(n33)
         );
  AOI22_X1 U75 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n11), .ZN(n29)
         );
  BUF_X1 U76 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U77 ( .A(sel), .Z(n1) );
  CLKBUF_X1 U78 ( .A(sel), .Z(n2) );
  INV_X1 U79 ( .A(n15), .ZN(n6) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_81 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  CLKBUF_X1 U1 ( .A(n3), .Z(n14) );
  CLKBUF_X1 U2 ( .A(n1), .Z(n7) );
  CLKBUF_X1 U3 ( .A(n1), .Z(n9) );
  BUF_X1 U4 ( .A(n3), .Z(n15) );
  INV_X1 U5 ( .A(n15), .ZN(n4) );
  INV_X1 U6 ( .A(n15), .ZN(n5) );
  INV_X1 U7 ( .A(n57), .ZN(N6) );
  AOI22_X1 U8 ( .A1(port0[4]), .A2(n6), .B1(port1[4]), .B2(n7), .ZN(n57) );
  INV_X1 U9 ( .A(n53), .ZN(N32) );
  AOI22_X1 U10 ( .A1(port0[30]), .A2(n6), .B1(port1[30]), .B2(n8), .ZN(n53) );
  INV_X1 U11 ( .A(n59), .ZN(N8) );
  AOI22_X1 U12 ( .A1(port0[6]), .A2(n6), .B1(port1[6]), .B2(n7), .ZN(n59) );
  INV_X1 U13 ( .A(n58), .ZN(N7) );
  AOI22_X1 U14 ( .A1(port0[5]), .A2(n6), .B1(port1[5]), .B2(n7), .ZN(n58) );
  INV_X1 U15 ( .A(n26), .ZN(N2) );
  AOI22_X1 U16 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n12), .ZN(n26) );
  INV_X1 U17 ( .A(n17), .ZN(N11) );
  AOI22_X1 U18 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n14), .ZN(n17) );
  INV_X1 U19 ( .A(n35), .ZN(N27) );
  AOI22_X1 U20 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n9), .ZN(n35) );
  INV_X1 U21 ( .A(n51), .ZN(N30) );
  AOI22_X1 U22 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n8), .ZN(n51) );
  INV_X1 U23 ( .A(n29), .ZN(N22) );
  AOI22_X1 U24 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n11), .ZN(n29)
         );
  INV_X1 U25 ( .A(n48), .ZN(N28) );
  AOI22_X1 U26 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n9), .ZN(n48) );
  INV_X1 U27 ( .A(n50), .ZN(N3) );
  AOI22_X1 U28 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n9), .ZN(n50) );
  INV_X1 U29 ( .A(n52), .ZN(N31) );
  AOI22_X1 U30 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n11), .ZN(n52)
         );
  INV_X1 U31 ( .A(n49), .ZN(N29) );
  AOI22_X1 U32 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n9), .ZN(n49) );
  INV_X1 U33 ( .A(n23), .ZN(N17) );
  AOI22_X1 U34 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n12), .ZN(n23)
         );
  INV_X1 U35 ( .A(n18), .ZN(N12) );
  AOI22_X1 U36 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n14), .ZN(n18)
         );
  INV_X1 U37 ( .A(n20), .ZN(N14) );
  AOI22_X1 U38 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n13), .ZN(n20)
         );
  INV_X1 U39 ( .A(n30), .ZN(N23) );
  AOI22_X1 U40 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n10), .ZN(n30)
         );
  INV_X1 U41 ( .A(n16), .ZN(N10) );
  AOI22_X1 U42 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n14), .ZN(n16) );
  INV_X1 U43 ( .A(n32), .ZN(N25) );
  AOI22_X1 U44 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n10), .ZN(n32)
         );
  INV_X1 U45 ( .A(n19), .ZN(N13) );
  AOI22_X1 U46 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n13), .ZN(n19)
         );
  INV_X1 U47 ( .A(n27), .ZN(N20) );
  AOI22_X1 U48 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n11), .ZN(n27)
         );
  INV_X1 U49 ( .A(n31), .ZN(N24) );
  AOI22_X1 U50 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n10), .ZN(n31)
         );
  INV_X1 U51 ( .A(n24), .ZN(N18) );
  AOI22_X1 U52 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n12), .ZN(n24)
         );
  INV_X1 U53 ( .A(n21), .ZN(N15) );
  AOI22_X1 U54 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n13), .ZN(n21)
         );
  INV_X1 U55 ( .A(n60), .ZN(N9) );
  AOI22_X1 U56 ( .A1(port0[7]), .A2(n6), .B1(n14), .B2(port1[7]), .ZN(n60) );
  INV_X1 U57 ( .A(n54), .ZN(N33) );
  AOI22_X1 U58 ( .A1(port0[31]), .A2(n6), .B1(port1[31]), .B2(n8), .ZN(n54) );
  INV_X1 U59 ( .A(n55), .ZN(N4) );
  AOI22_X1 U60 ( .A1(port0[2]), .A2(n6), .B1(port1[2]), .B2(n8), .ZN(n55) );
  INV_X1 U61 ( .A(n56), .ZN(N5) );
  AOI22_X1 U62 ( .A1(port0[3]), .A2(n6), .B1(port1[3]), .B2(n7), .ZN(n56) );
  BUF_X1 U63 ( .A(n1), .Z(n8) );
  BUF_X1 U64 ( .A(n2), .Z(n12) );
  BUF_X1 U65 ( .A(n2), .Z(n11) );
  BUF_X1 U66 ( .A(n2), .Z(n10) );
  BUF_X1 U67 ( .A(n3), .Z(n13) );
  INV_X1 U68 ( .A(n22), .ZN(N16) );
  AOI22_X1 U69 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n13), .ZN(n22)
         );
  INV_X1 U70 ( .A(n25), .ZN(N19) );
  AOI22_X1 U71 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n12), .ZN(n25)
         );
  INV_X1 U72 ( .A(n28), .ZN(N21) );
  AOI22_X1 U73 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n11), .ZN(n28)
         );
  INV_X1 U74 ( .A(n33), .ZN(N26) );
  AOI22_X1 U75 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n10), .ZN(n33)
         );
  BUF_X1 U76 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U77 ( .A(sel), .Z(n1) );
  CLKBUF_X1 U78 ( .A(sel), .Z(n2) );
  INV_X1 U79 ( .A(n15), .ZN(n6) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_80 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n40, n41, n45, net132913, net132909, net132907,
         net132903, net132901, net132893, net132919, net149162, net169428,
         net169505, net169633, net169648, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23,
         n24, n25, n26, n27, n28, n29, n30, n31, n32;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  BUF_X2 U1 ( .A(net149162), .Z(net132907) );
  CLKBUF_X3 U2 ( .A(net132919), .Z(net132913) );
  CLKBUF_X1 U3 ( .A(sel), .Z(net132919) );
  CLKBUF_X1 U4 ( .A(net132919), .Z(net132909) );
  CLKBUF_X1 U5 ( .A(net132919), .Z(net132903) );
  BUF_X1 U6 ( .A(n4), .Z(net149162) );
  INV_X1 U7 ( .A(net132913), .ZN(n1) );
  INV_X1 U8 ( .A(net132909), .ZN(net132893) );
  BUF_X1 U9 ( .A(sel), .Z(n4) );
  BUF_X1 U10 ( .A(net149162), .Z(net132901) );
  AOI22_X1 U11 ( .A1(port0[0]), .A2(net169633), .B1(port1[0]), .B2(net132913), 
        .ZN(n2) );
  INV_X1 U12 ( .A(n2), .ZN(N2) );
  INV_X1 U13 ( .A(net132909), .ZN(n3) );
  AOI22_X1 U14 ( .A1(port0[1]), .A2(n3), .B1(port1[1]), .B2(net132903), .ZN(
        n45) );
  AOI22_X1 U15 ( .A1(port0[31]), .A2(n1), .B1(port1[31]), .B2(net132901), .ZN(
        n41) );
  AOI22_X1 U16 ( .A1(port0[2]), .A2(n3), .B1(port1[2]), .B2(net132901), .ZN(
        n40) );
  CLKBUF_X1 U17 ( .A(sel), .Z(net169648) );
  INV_X1 U18 ( .A(sel), .ZN(net169428) );
  INV_X1 U19 ( .A(net149162), .ZN(net169633) );
  INV_X1 U20 ( .A(net132913), .ZN(net169505) );
  INV_X1 U21 ( .A(n27), .ZN(N32) );
  INV_X1 U22 ( .A(n41), .ZN(N33) );
  INV_X1 U23 ( .A(n23), .ZN(N28) );
  INV_X1 U24 ( .A(n19), .ZN(N24) );
  INV_X1 U25 ( .A(n18), .ZN(N23) );
  INV_X1 U26 ( .A(n26), .ZN(N31) );
  INV_X1 U27 ( .A(n24), .ZN(N29) );
  INV_X1 U28 ( .A(n25), .ZN(N30) );
  INV_X1 U29 ( .A(n22), .ZN(N27) );
  INV_X1 U30 ( .A(n20), .ZN(N25) );
  INV_X1 U31 ( .A(n16), .ZN(N21) );
  INV_X1 U32 ( .A(n21), .ZN(N26) );
  INV_X1 U33 ( .A(n17), .ZN(N22) );
  INV_X1 U34 ( .A(n15), .ZN(N20) );
  INV_X1 U35 ( .A(n14), .ZN(N19) );
  INV_X1 U36 ( .A(n13), .ZN(N18) );
  INV_X1 U37 ( .A(n29), .ZN(N6) );
  AOI22_X1 U38 ( .A1(port0[26]), .A2(net169505), .B1(port1[26]), .B2(net132913), .ZN(n23) );
  AOI22_X1 U39 ( .A1(port0[21]), .A2(net169505), .B1(port1[21]), .B2(net132907), .ZN(n18) );
  AOI22_X1 U40 ( .A1(port0[29]), .A2(n1), .B1(port1[29]), .B2(net132907), .ZN(
        n26) );
  AOI22_X1 U41 ( .A1(port0[25]), .A2(n1), .B1(port1[25]), .B2(net132903), .ZN(
        n22) );
  AOI22_X1 U42 ( .A1(port0[28]), .A2(net169505), .B1(port1[28]), .B2(net132901), .ZN(n25) );
  AOI22_X1 U43 ( .A1(port0[20]), .A2(net132893), .B1(port1[20]), .B2(net132907), .ZN(n17) );
  AOI22_X1 U44 ( .A1(port0[24]), .A2(net132893), .B1(port1[24]), .B2(net132907), .ZN(n21) );
  INV_X1 U45 ( .A(n40), .ZN(N4) );
  INV_X1 U46 ( .A(n45), .ZN(N3) );
  INV_X1 U47 ( .A(n28), .ZN(N5) );
  INV_X1 U48 ( .A(n30), .ZN(N7) );
  INV_X1 U49 ( .A(n31), .ZN(N8) );
  INV_X1 U50 ( .A(n9), .ZN(N14) );
  INV_X1 U51 ( .A(n8), .ZN(N13) );
  INV_X1 U52 ( .A(n11), .ZN(N16) );
  INV_X1 U53 ( .A(n5), .ZN(N10) );
  INV_X1 U54 ( .A(n6), .ZN(N11) );
  INV_X1 U55 ( .A(n10), .ZN(N15) );
  INV_X1 U56 ( .A(n7), .ZN(N12) );
  AOI22_X1 U57 ( .A1(port0[22]), .A2(n1), .B1(port1[22]), .B2(net132907), .ZN(
        n19) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(net169505), .B1(port1[19]), .B2(net132907), .ZN(n16) );
  AOI22_X1 U59 ( .A1(port0[27]), .A2(net169633), .B1(port1[27]), .B2(net132913), .ZN(n24) );
  AOI22_X1 U60 ( .A1(port0[23]), .A2(n1), .B1(port1[23]), .B2(net132907), .ZN(
        n20) );
  AOI22_X1 U61 ( .A1(port0[16]), .A2(net169505), .B1(port1[16]), .B2(net132903), .ZN(n13) );
  AOI22_X1 U62 ( .A1(port0[18]), .A2(n1), .B1(port1[18]), .B2(net132907), .ZN(
        n15) );
  AOI22_X1 U63 ( .A1(port0[17]), .A2(net132893), .B1(port1[17]), .B2(net132913), .ZN(n14) );
  AOI22_X1 U64 ( .A1(port0[11]), .A2(net169505), .B1(port1[11]), .B2(net132903), .ZN(n8) );
  AOI22_X1 U65 ( .A1(port0[13]), .A2(net132893), .B1(port1[13]), .B2(net132903), .ZN(n10) );
  AOI22_X1 U66 ( .A1(port0[12]), .A2(net169505), .B1(port1[12]), .B2(net132913), .ZN(n9) );
  AOI22_X1 U67 ( .A1(port0[14]), .A2(net132893), .B1(port1[14]), .B2(net132913), .ZN(n11) );
  AOI22_X1 U68 ( .A1(port0[8]), .A2(net169633), .B1(port1[8]), .B2(net132913), 
        .ZN(n5) );
  AOI22_X1 U69 ( .A1(port0[10]), .A2(n1), .B1(port1[10]), .B2(net132913), .ZN(
        n7) );
  AOI22_X1 U70 ( .A1(port0[9]), .A2(net132893), .B1(port1[9]), .B2(net132903), 
        .ZN(n6) );
  INV_X1 U71 ( .A(n12), .ZN(N17) );
  AOI22_X1 U72 ( .A1(net169428), .A2(port0[15]), .B1(n4), .B2(port1[15]), .ZN(
        n12) );
  AOI22_X1 U73 ( .A1(port0[30]), .A2(net169505), .B1(port1[30]), .B2(net132901), .ZN(n27) );
  AOI22_X1 U74 ( .A1(port0[5]), .A2(net132893), .B1(port1[5]), .B2(net132907), 
        .ZN(n30) );
  AOI22_X1 U75 ( .A1(port0[6]), .A2(n1), .B1(port1[6]), .B2(net132907), .ZN(
        n31) );
  AOI22_X1 U76 ( .A1(port0[4]), .A2(net169633), .B1(port1[4]), .B2(net132907), 
        .ZN(n29) );
  AOI22_X1 U77 ( .A1(port0[3]), .A2(net132893), .B1(port1[3]), .B2(net132907), 
        .ZN(n28) );
  AOI22_X1 U78 ( .A1(net169428), .A2(port0[7]), .B1(net169648), .B2(port1[7]), 
        .ZN(n32) );
  INV_X1 U79 ( .A(n32), .ZN(N9) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_51 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n25), .ZN(N2) );
  INV_X1 U2 ( .A(n55), .ZN(N6) );
  INV_X1 U3 ( .A(n54), .ZN(N5) );
  INV_X1 U4 ( .A(n53), .ZN(N4) );
  INV_X1 U5 ( .A(n48), .ZN(N3) );
  INV_X1 U6 ( .A(n14), .ZN(n4) );
  INV_X1 U7 ( .A(n58), .ZN(N9) );
  INV_X1 U8 ( .A(n56), .ZN(N7) );
  INV_X1 U9 ( .A(n57), .ZN(N8) );
  INV_X1 U10 ( .A(n17), .ZN(N12) );
  INV_X1 U11 ( .A(n52), .ZN(N33) );
  INV_X1 U12 ( .A(n51), .ZN(N32) );
  INV_X1 U13 ( .A(n26), .ZN(N20) );
  INV_X1 U14 ( .A(n20), .ZN(N15) );
  INV_X1 U15 ( .A(n19), .ZN(N14) );
  INV_X1 U16 ( .A(n21), .ZN(N16) );
  INV_X1 U17 ( .A(n18), .ZN(N13) );
  INV_X1 U18 ( .A(n27), .ZN(N21) );
  INV_X1 U19 ( .A(n28), .ZN(N22) );
  INV_X1 U20 ( .A(n29), .ZN(N23) );
  INV_X1 U21 ( .A(n30), .ZN(N24) );
  INV_X1 U22 ( .A(n31), .ZN(N25) );
  INV_X1 U23 ( .A(n32), .ZN(N26) );
  INV_X1 U24 ( .A(n33), .ZN(N27) );
  INV_X1 U25 ( .A(n35), .ZN(N28) );
  INV_X1 U26 ( .A(n47), .ZN(N29) );
  INV_X1 U27 ( .A(n49), .ZN(N30) );
  INV_X1 U28 ( .A(n50), .ZN(N31) );
  INV_X1 U29 ( .A(n16), .ZN(N11) );
  INV_X1 U30 ( .A(n15), .ZN(N10) );
  INV_X1 U31 ( .A(n24), .ZN(N19) );
  INV_X1 U32 ( .A(n22), .ZN(N17) );
  INV_X1 U33 ( .A(n23), .ZN(N18) );
  INV_X1 U34 ( .A(n14), .ZN(n5) );
  AOI22_X1 U35 ( .A1(port0[4]), .A2(n5), .B1(port1[4]), .B2(n6), .ZN(n55) );
  AOI22_X1 U36 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  AOI22_X1 U37 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  AOI22_X1 U38 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  AOI22_X1 U39 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(n7), .ZN(n53) );
  AOI22_X1 U40 ( .A1(port0[7]), .A2(n5), .B1(n13), .B2(port1[7]), .ZN(n58) );
  AOI22_X1 U41 ( .A1(port0[6]), .A2(n5), .B1(port1[6]), .B2(n6), .ZN(n57) );
  AOI22_X1 U42 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  AOI22_X1 U43 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  AOI22_X1 U45 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  AOI22_X1 U46 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  AOI22_X1 U47 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  AOI22_X1 U48 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  AOI22_X1 U49 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  BUF_X1 U50 ( .A(n2), .Z(n11) );
  BUF_X1 U51 ( .A(n3), .Z(n14) );
  AOI22_X1 U52 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  AOI22_X1 U53 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n7), .ZN(n52) );
  AOI22_X1 U54 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n7), .ZN(n51) );
  AOI22_X1 U55 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  AOI22_X1 U56 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  AOI22_X1 U57 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  AOI22_X1 U58 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  AOI22_X1 U59 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  AOI22_X1 U60 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  AOI22_X1 U61 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  AOI22_X1 U62 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  AOI22_X1 U63 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  AOI22_X1 U64 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  AOI22_X1 U65 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  AOI22_X1 U66 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  AOI22_X1 U67 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  AOI22_X1 U68 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  BUF_X1 U69 ( .A(n1), .Z(n6) );
  BUF_X1 U70 ( .A(n1), .Z(n8) );
  BUF_X1 U71 ( .A(n1), .Z(n7) );
  BUF_X1 U72 ( .A(n3), .Z(n13) );
  BUF_X1 U73 ( .A(n3), .Z(n12) );
  BUF_X1 U74 ( .A(n2), .Z(n10) );
  BUF_X1 U75 ( .A(n2), .Z(n9) );
  BUF_X1 U76 ( .A(sel), .Z(n3) );
  BUF_X1 U77 ( .A(sel), .Z(n2) );
  BUF_X1 U78 ( .A(sel), .Z(n1) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_50 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n25), .ZN(N2) );
  INV_X1 U2 ( .A(n55), .ZN(N6) );
  INV_X1 U3 ( .A(n54), .ZN(N5) );
  INV_X1 U4 ( .A(n53), .ZN(N4) );
  INV_X1 U5 ( .A(n48), .ZN(N3) );
  INV_X1 U6 ( .A(n14), .ZN(n4) );
  INV_X1 U7 ( .A(n58), .ZN(N9) );
  INV_X1 U8 ( .A(n56), .ZN(N7) );
  INV_X1 U9 ( .A(n57), .ZN(N8) );
  INV_X1 U10 ( .A(n17), .ZN(N12) );
  INV_X1 U11 ( .A(n52), .ZN(N33) );
  INV_X1 U12 ( .A(n51), .ZN(N32) );
  INV_X1 U13 ( .A(n26), .ZN(N20) );
  INV_X1 U14 ( .A(n20), .ZN(N15) );
  INV_X1 U15 ( .A(n19), .ZN(N14) );
  INV_X1 U16 ( .A(n21), .ZN(N16) );
  INV_X1 U17 ( .A(n18), .ZN(N13) );
  INV_X1 U18 ( .A(n27), .ZN(N21) );
  INV_X1 U19 ( .A(n28), .ZN(N22) );
  INV_X1 U20 ( .A(n29), .ZN(N23) );
  INV_X1 U21 ( .A(n30), .ZN(N24) );
  INV_X1 U22 ( .A(n31), .ZN(N25) );
  INV_X1 U23 ( .A(n32), .ZN(N26) );
  INV_X1 U24 ( .A(n33), .ZN(N27) );
  INV_X1 U25 ( .A(n35), .ZN(N28) );
  INV_X1 U26 ( .A(n47), .ZN(N29) );
  INV_X1 U27 ( .A(n49), .ZN(N30) );
  INV_X1 U28 ( .A(n50), .ZN(N31) );
  INV_X1 U29 ( .A(n16), .ZN(N11) );
  INV_X1 U30 ( .A(n15), .ZN(N10) );
  INV_X1 U31 ( .A(n24), .ZN(N19) );
  INV_X1 U32 ( .A(n22), .ZN(N17) );
  INV_X1 U33 ( .A(n23), .ZN(N18) );
  INV_X1 U34 ( .A(n14), .ZN(n5) );
  AOI22_X1 U35 ( .A1(port0[4]), .A2(n5), .B1(port1[4]), .B2(n6), .ZN(n55) );
  AOI22_X1 U36 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  AOI22_X1 U37 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(n7), .ZN(n53) );
  AOI22_X1 U38 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  AOI22_X1 U39 ( .A1(port0[7]), .A2(n5), .B1(n13), .B2(port1[7]), .ZN(n58) );
  AOI22_X1 U40 ( .A1(port0[6]), .A2(n5), .B1(port1[6]), .B2(n6), .ZN(n57) );
  AOI22_X1 U41 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  AOI22_X1 U42 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  AOI22_X1 U43 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  AOI22_X1 U45 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  AOI22_X1 U46 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  AOI22_X1 U47 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  AOI22_X1 U48 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  AOI22_X1 U49 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  BUF_X1 U50 ( .A(n3), .Z(n14) );
  BUF_X1 U51 ( .A(n2), .Z(n11) );
  AOI22_X1 U52 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  AOI22_X1 U53 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n7), .ZN(n52) );
  AOI22_X1 U54 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n7), .ZN(n51) );
  AOI22_X1 U55 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  AOI22_X1 U56 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  AOI22_X1 U57 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  AOI22_X1 U58 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  AOI22_X1 U59 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  AOI22_X1 U60 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  AOI22_X1 U61 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  AOI22_X1 U62 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  AOI22_X1 U63 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  AOI22_X1 U64 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  AOI22_X1 U65 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  AOI22_X1 U66 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  AOI22_X1 U67 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  BUF_X1 U68 ( .A(n1), .Z(n6) );
  BUF_X1 U69 ( .A(n1), .Z(n8) );
  BUF_X1 U70 ( .A(n1), .Z(n7) );
  BUF_X1 U71 ( .A(n3), .Z(n13) );
  BUF_X1 U72 ( .A(n3), .Z(n12) );
  BUF_X1 U73 ( .A(n2), .Z(n10) );
  BUF_X1 U74 ( .A(n2), .Z(n9) );
  BUF_X1 U75 ( .A(sel), .Z(n3) );
  BUF_X1 U76 ( .A(sel), .Z(n2) );
  BUF_X1 U77 ( .A(sel), .Z(n1) );
  AOI22_X1 U78 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_49 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  AOI22_X1 U1 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  INV_X1 U2 ( .A(n55), .ZN(N6) );
  AOI22_X1 U3 ( .A1(port0[4]), .A2(n5), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U4 ( .A(n54), .ZN(N5) );
  AOI22_X1 U5 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U6 ( .A(n53), .ZN(N4) );
  AOI22_X1 U7 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U8 ( .A(n48), .ZN(N3) );
  AOI22_X1 U9 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  INV_X1 U10 ( .A(n14), .ZN(n4) );
  INV_X1 U11 ( .A(n58), .ZN(N9) );
  AOI22_X1 U12 ( .A1(port0[7]), .A2(n5), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U13 ( .A(n56), .ZN(N7) );
  AOI22_X1 U14 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U15 ( .A(n57), .ZN(N8) );
  AOI22_X1 U16 ( .A1(port0[6]), .A2(n5), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U17 ( .A(n17), .ZN(N12) );
  AOI22_X1 U18 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U19 ( .A(n52), .ZN(N33) );
  AOI22_X1 U20 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n7), .ZN(n52) );
  INV_X1 U21 ( .A(n51), .ZN(N32) );
  AOI22_X1 U22 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n7), .ZN(n51) );
  INV_X1 U23 ( .A(n26), .ZN(N20) );
  AOI22_X1 U24 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  INV_X1 U25 ( .A(n20), .ZN(N15) );
  AOI22_X1 U26 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U27 ( .A(n19), .ZN(N14) );
  AOI22_X1 U28 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U29 ( .A(n21), .ZN(N16) );
  AOI22_X1 U30 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U31 ( .A(n18), .ZN(N13) );
  AOI22_X1 U32 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U33 ( .A(n27), .ZN(N21) );
  AOI22_X1 U34 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  INV_X1 U35 ( .A(n28), .ZN(N22) );
  AOI22_X1 U36 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U37 ( .A(n29), .ZN(N23) );
  AOI22_X1 U38 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  INV_X1 U39 ( .A(n30), .ZN(N24) );
  AOI22_X1 U40 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  INV_X1 U41 ( .A(n31), .ZN(N25) );
  AOI22_X1 U42 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  INV_X1 U43 ( .A(n32), .ZN(N26) );
  AOI22_X1 U44 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U45 ( .A(n33), .ZN(N27) );
  AOI22_X1 U46 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  INV_X1 U47 ( .A(n35), .ZN(N28) );
  AOI22_X1 U48 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  INV_X1 U49 ( .A(n47), .ZN(N29) );
  AOI22_X1 U50 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  INV_X1 U51 ( .A(n49), .ZN(N30) );
  AOI22_X1 U52 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U53 ( .A(n50), .ZN(N31) );
  AOI22_X1 U54 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  INV_X1 U55 ( .A(n16), .ZN(N11) );
  AOI22_X1 U56 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U57 ( .A(n15), .ZN(N10) );
  AOI22_X1 U58 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U59 ( .A(n24), .ZN(N19) );
  AOI22_X1 U60 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U61 ( .A(n22), .ZN(N17) );
  AOI22_X1 U62 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  INV_X1 U63 ( .A(n23), .ZN(N18) );
  AOI22_X1 U64 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  BUF_X1 U65 ( .A(n3), .Z(n14) );
  BUF_X1 U66 ( .A(n2), .Z(n11) );
  BUF_X1 U67 ( .A(n1), .Z(n8) );
  BUF_X1 U68 ( .A(n1), .Z(n7) );
  BUF_X1 U69 ( .A(n1), .Z(n6) );
  BUF_X1 U70 ( .A(n3), .Z(n13) );
  BUF_X1 U71 ( .A(n3), .Z(n12) );
  BUF_X1 U72 ( .A(n2), .Z(n10) );
  BUF_X1 U73 ( .A(n2), .Z(n9) );
  BUF_X1 U74 ( .A(sel), .Z(n3) );
  BUF_X1 U75 ( .A(sel), .Z(n2) );
  BUF_X1 U76 ( .A(sel), .Z(n1) );
  INV_X1 U77 ( .A(n25), .ZN(N2) );
  INV_X1 U78 ( .A(n14), .ZN(n5) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_20 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  INV_X1 U3 ( .A(n53), .ZN(N4) );
  AOI22_X1 U4 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U5 ( .A(n54), .ZN(N5) );
  AOI22_X1 U6 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U7 ( .A(n55), .ZN(N6) );
  AOI22_X1 U8 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U9 ( .A(n56), .ZN(N7) );
  AOI22_X1 U10 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U11 ( .A(n57), .ZN(N8) );
  AOI22_X1 U12 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U13 ( .A(n58), .ZN(N9) );
  AOI22_X1 U14 ( .A1(port0[7]), .A2(n5), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U15 ( .A(n51), .ZN(N32) );
  AOI22_X1 U16 ( .A1(port0[30]), .A2(n4), .B1(port1[30]), .B2(n7), .ZN(n51) );
  INV_X1 U17 ( .A(n52), .ZN(N33) );
  AOI22_X1 U18 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n7), .ZN(n52) );
  INV_X1 U19 ( .A(n25), .ZN(N2) );
  AOI22_X1 U20 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  INV_X1 U21 ( .A(n48), .ZN(N3) );
  AOI22_X1 U22 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  INV_X1 U23 ( .A(n18), .ZN(N13) );
  AOI22_X1 U24 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U25 ( .A(n19), .ZN(N14) );
  AOI22_X1 U26 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U27 ( .A(n20), .ZN(N15) );
  AOI22_X1 U28 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U29 ( .A(n21), .ZN(N16) );
  AOI22_X1 U30 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U31 ( .A(n22), .ZN(N17) );
  AOI22_X1 U32 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  INV_X1 U33 ( .A(n23), .ZN(N18) );
  AOI22_X1 U34 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  INV_X1 U35 ( .A(n24), .ZN(N19) );
  AOI22_X1 U36 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U37 ( .A(n26), .ZN(N20) );
  AOI22_X1 U38 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  INV_X1 U39 ( .A(n27), .ZN(N21) );
  AOI22_X1 U40 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  INV_X1 U41 ( .A(n28), .ZN(N22) );
  AOI22_X1 U42 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U43 ( .A(n29), .ZN(N23) );
  AOI22_X1 U44 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  INV_X1 U45 ( .A(n30), .ZN(N24) );
  AOI22_X1 U46 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  INV_X1 U47 ( .A(n31), .ZN(N25) );
  AOI22_X1 U48 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  INV_X1 U49 ( .A(n32), .ZN(N26) );
  AOI22_X1 U50 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U51 ( .A(n33), .ZN(N27) );
  AOI22_X1 U52 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  INV_X1 U53 ( .A(n35), .ZN(N28) );
  AOI22_X1 U54 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  INV_X1 U55 ( .A(n47), .ZN(N29) );
  AOI22_X1 U56 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  INV_X1 U57 ( .A(n49), .ZN(N30) );
  AOI22_X1 U58 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U59 ( .A(n50), .ZN(N31) );
  AOI22_X1 U60 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  INV_X1 U61 ( .A(n15), .ZN(N10) );
  AOI22_X1 U62 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U63 ( .A(n16), .ZN(N11) );
  AOI22_X1 U64 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U65 ( .A(n17), .ZN(N12) );
  AOI22_X1 U66 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  BUF_X1 U67 ( .A(n1), .Z(n6) );
  BUF_X1 U68 ( .A(n3), .Z(n12) );
  BUF_X1 U69 ( .A(n2), .Z(n11) );
  BUF_X1 U70 ( .A(n2), .Z(n9) );
  BUF_X1 U71 ( .A(n1), .Z(n8) );
  BUF_X1 U72 ( .A(n2), .Z(n10) );
  BUF_X1 U73 ( .A(n1), .Z(n7) );
  BUF_X1 U74 ( .A(n3), .Z(n14) );
  BUF_X1 U75 ( .A(n3), .Z(n13) );
  BUF_X1 U76 ( .A(sel), .Z(n3) );
  BUF_X1 U77 ( .A(sel), .Z(n2) );
  BUF_X1 U78 ( .A(sel), .Z(n1) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_19 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  INV_X1 U3 ( .A(n58), .ZN(N9) );
  AOI22_X1 U4 ( .A1(port0[7]), .A2(n4), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U5 ( .A(n53), .ZN(N4) );
  AOI22_X1 U6 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U7 ( .A(n54), .ZN(N5) );
  AOI22_X1 U8 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U9 ( .A(n55), .ZN(N6) );
  AOI22_X1 U10 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U11 ( .A(n56), .ZN(N7) );
  AOI22_X1 U12 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U13 ( .A(n57), .ZN(N8) );
  AOI22_X1 U14 ( .A1(port0[6]), .A2(n5), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U15 ( .A(n51), .ZN(N32) );
  AOI22_X1 U16 ( .A1(port0[30]), .A2(n4), .B1(port1[30]), .B2(n7), .ZN(n51) );
  INV_X1 U17 ( .A(n52), .ZN(N33) );
  AOI22_X1 U18 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n7), .ZN(n52) );
  INV_X1 U19 ( .A(n25), .ZN(N2) );
  AOI22_X1 U20 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  INV_X1 U21 ( .A(n48), .ZN(N3) );
  AOI22_X1 U22 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  INV_X1 U23 ( .A(n18), .ZN(N13) );
  AOI22_X1 U24 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U25 ( .A(n19), .ZN(N14) );
  AOI22_X1 U26 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U27 ( .A(n20), .ZN(N15) );
  AOI22_X1 U28 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U29 ( .A(n21), .ZN(N16) );
  AOI22_X1 U30 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U31 ( .A(n22), .ZN(N17) );
  AOI22_X1 U32 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  INV_X1 U33 ( .A(n23), .ZN(N18) );
  AOI22_X1 U34 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  INV_X1 U35 ( .A(n24), .ZN(N19) );
  AOI22_X1 U36 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U37 ( .A(n26), .ZN(N20) );
  AOI22_X1 U38 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  INV_X1 U39 ( .A(n27), .ZN(N21) );
  AOI22_X1 U40 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  INV_X1 U41 ( .A(n28), .ZN(N22) );
  AOI22_X1 U42 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U43 ( .A(n29), .ZN(N23) );
  AOI22_X1 U44 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  INV_X1 U45 ( .A(n30), .ZN(N24) );
  AOI22_X1 U46 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  INV_X1 U47 ( .A(n31), .ZN(N25) );
  AOI22_X1 U48 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  INV_X1 U49 ( .A(n32), .ZN(N26) );
  AOI22_X1 U50 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U51 ( .A(n33), .ZN(N27) );
  AOI22_X1 U52 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  INV_X1 U53 ( .A(n35), .ZN(N28) );
  AOI22_X1 U54 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  INV_X1 U55 ( .A(n47), .ZN(N29) );
  AOI22_X1 U56 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  INV_X1 U57 ( .A(n49), .ZN(N30) );
  AOI22_X1 U58 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U59 ( .A(n50), .ZN(N31) );
  AOI22_X1 U60 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  INV_X1 U61 ( .A(n15), .ZN(N10) );
  AOI22_X1 U62 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U63 ( .A(n16), .ZN(N11) );
  AOI22_X1 U64 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U65 ( .A(n17), .ZN(N12) );
  AOI22_X1 U66 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  BUF_X1 U67 ( .A(n1), .Z(n6) );
  BUF_X1 U68 ( .A(n3), .Z(n12) );
  BUF_X1 U69 ( .A(n2), .Z(n11) );
  BUF_X1 U70 ( .A(n2), .Z(n9) );
  BUF_X1 U71 ( .A(n1), .Z(n8) );
  BUF_X1 U72 ( .A(n2), .Z(n10) );
  BUF_X1 U73 ( .A(n1), .Z(n7) );
  BUF_X1 U74 ( .A(n3), .Z(n14) );
  BUF_X1 U75 ( .A(n3), .Z(n13) );
  BUF_X1 U76 ( .A(sel), .Z(n3) );
  BUF_X1 U77 ( .A(sel), .Z(n2) );
  BUF_X1 U78 ( .A(sel), .Z(n1) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_18 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  BUF_X1 U3 ( .A(n1), .Z(n6) );
  BUF_X1 U4 ( .A(n3), .Z(n12) );
  BUF_X1 U5 ( .A(n2), .Z(n11) );
  BUF_X1 U6 ( .A(n2), .Z(n9) );
  BUF_X1 U7 ( .A(n1), .Z(n8) );
  BUF_X1 U8 ( .A(n2), .Z(n10) );
  BUF_X1 U9 ( .A(n1), .Z(n7) );
  BUF_X1 U10 ( .A(n3), .Z(n14) );
  BUF_X1 U11 ( .A(n3), .Z(n13) );
  BUF_X1 U12 ( .A(sel), .Z(n3) );
  BUF_X1 U13 ( .A(sel), .Z(n2) );
  BUF_X1 U14 ( .A(sel), .Z(n1) );
  INV_X1 U15 ( .A(n25), .ZN(N2) );
  AOI22_X1 U16 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  INV_X1 U17 ( .A(n48), .ZN(N3) );
  AOI22_X1 U18 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  INV_X1 U19 ( .A(n33), .ZN(N27) );
  AOI22_X1 U20 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  INV_X1 U21 ( .A(n35), .ZN(N28) );
  AOI22_X1 U22 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  INV_X1 U23 ( .A(n47), .ZN(N29) );
  AOI22_X1 U24 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  INV_X1 U25 ( .A(n49), .ZN(N30) );
  AOI22_X1 U26 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U27 ( .A(n50), .ZN(N31) );
  AOI22_X1 U28 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  INV_X1 U29 ( .A(n51), .ZN(N32) );
  AOI22_X1 U30 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n7), .ZN(n51) );
  INV_X1 U31 ( .A(n53), .ZN(N4) );
  AOI22_X1 U32 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U33 ( .A(n54), .ZN(N5) );
  AOI22_X1 U34 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U35 ( .A(n55), .ZN(N6) );
  AOI22_X1 U36 ( .A1(port0[4]), .A2(n5), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U37 ( .A(n56), .ZN(N7) );
  AOI22_X1 U38 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U39 ( .A(n57), .ZN(N8) );
  AOI22_X1 U40 ( .A1(port0[6]), .A2(n5), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U41 ( .A(n58), .ZN(N9) );
  AOI22_X1 U42 ( .A1(port0[7]), .A2(n4), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U43 ( .A(n15), .ZN(N10) );
  AOI22_X1 U44 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U45 ( .A(n16), .ZN(N11) );
  AOI22_X1 U46 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U47 ( .A(n17), .ZN(N12) );
  AOI22_X1 U48 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U49 ( .A(n18), .ZN(N13) );
  AOI22_X1 U50 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U51 ( .A(n19), .ZN(N14) );
  AOI22_X1 U52 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U53 ( .A(n20), .ZN(N15) );
  AOI22_X1 U54 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U55 ( .A(n21), .ZN(N16) );
  AOI22_X1 U56 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U57 ( .A(n22), .ZN(N17) );
  AOI22_X1 U58 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  INV_X1 U59 ( .A(n23), .ZN(N18) );
  AOI22_X1 U60 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  INV_X1 U61 ( .A(n24), .ZN(N19) );
  AOI22_X1 U62 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U63 ( .A(n26), .ZN(N20) );
  AOI22_X1 U64 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  INV_X1 U65 ( .A(n27), .ZN(N21) );
  AOI22_X1 U66 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  INV_X1 U67 ( .A(n28), .ZN(N22) );
  AOI22_X1 U68 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U69 ( .A(n29), .ZN(N23) );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  INV_X1 U71 ( .A(n30), .ZN(N24) );
  AOI22_X1 U72 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  INV_X1 U73 ( .A(n31), .ZN(N25) );
  AOI22_X1 U74 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  INV_X1 U75 ( .A(n32), .ZN(N26) );
  AOI22_X1 U76 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U77 ( .A(n52), .ZN(N33) );
  AOI22_X1 U78 ( .A1(port0[31]), .A2(n4), .B1(port1[31]), .B2(n7), .ZN(n52) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_17 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n5) );
  INV_X1 U2 ( .A(n14), .ZN(n4) );
  BUF_X1 U3 ( .A(n1), .Z(n8) );
  BUF_X1 U4 ( .A(n1), .Z(n7) );
  BUF_X1 U5 ( .A(n1), .Z(n6) );
  BUF_X1 U6 ( .A(n3), .Z(n14) );
  BUF_X1 U7 ( .A(n3), .Z(n13) );
  BUF_X1 U8 ( .A(n2), .Z(n11) );
  BUF_X1 U9 ( .A(n3), .Z(n12) );
  BUF_X1 U10 ( .A(n2), .Z(n10) );
  BUF_X1 U11 ( .A(n2), .Z(n9) );
  INV_X1 U12 ( .A(n28), .ZN(N22) );
  AOI22_X1 U13 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U14 ( .A(n29), .ZN(N23) );
  AOI22_X1 U15 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  INV_X1 U16 ( .A(n30), .ZN(N24) );
  AOI22_X1 U17 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  INV_X1 U18 ( .A(n31), .ZN(N25) );
  AOI22_X1 U19 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  INV_X1 U20 ( .A(n32), .ZN(N26) );
  AOI22_X1 U21 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U22 ( .A(n33), .ZN(N27) );
  AOI22_X1 U23 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  INV_X1 U24 ( .A(n35), .ZN(N28) );
  AOI22_X1 U25 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  INV_X1 U26 ( .A(n47), .ZN(N29) );
  AOI22_X1 U27 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  INV_X1 U28 ( .A(n26), .ZN(N20) );
  AOI22_X1 U29 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  INV_X1 U30 ( .A(n24), .ZN(N19) );
  AOI22_X1 U31 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U32 ( .A(n23), .ZN(N18) );
  AOI22_X1 U33 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  INV_X1 U34 ( .A(n27), .ZN(N21) );
  AOI22_X1 U35 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  INV_X1 U36 ( .A(n52), .ZN(N33) );
  AOI22_X1 U37 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n7), .ZN(n52) );
  INV_X1 U38 ( .A(n49), .ZN(N30) );
  AOI22_X1 U39 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U40 ( .A(n50), .ZN(N31) );
  AOI22_X1 U41 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  INV_X1 U42 ( .A(n51), .ZN(N32) );
  AOI22_X1 U43 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n7), .ZN(n51) );
  BUF_X1 U44 ( .A(sel), .Z(n3) );
  BUF_X1 U45 ( .A(sel), .Z(n2) );
  BUF_X1 U46 ( .A(sel), .Z(n1) );
  INV_X1 U47 ( .A(n55), .ZN(N6) );
  AOI22_X1 U48 ( .A1(port0[4]), .A2(n5), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U49 ( .A(n54), .ZN(N5) );
  AOI22_X1 U50 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U51 ( .A(n53), .ZN(N4) );
  AOI22_X1 U52 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U53 ( .A(n25), .ZN(N2) );
  INV_X1 U54 ( .A(n48), .ZN(N3) );
  AOI22_X1 U55 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  INV_X1 U56 ( .A(n22), .ZN(N17) );
  AOI22_X1 U57 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  INV_X1 U58 ( .A(n56), .ZN(N7) );
  AOI22_X1 U59 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U60 ( .A(n58), .ZN(N9) );
  AOI22_X1 U61 ( .A1(port0[7]), .A2(n5), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U62 ( .A(n57), .ZN(N8) );
  AOI22_X1 U63 ( .A1(port0[6]), .A2(n5), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U64 ( .A(n20), .ZN(N15) );
  AOI22_X1 U65 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U66 ( .A(n19), .ZN(N14) );
  AOI22_X1 U67 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U68 ( .A(n21), .ZN(N16) );
  AOI22_X1 U69 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U70 ( .A(n18), .ZN(N13) );
  AOI22_X1 U71 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U72 ( .A(n17), .ZN(N12) );
  AOI22_X1 U73 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U74 ( .A(n16), .ZN(N11) );
  AOI22_X1 U75 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U76 ( .A(n15), .ZN(N10) );
  AOI22_X1 U77 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  AOI22_X1 U78 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_16 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  BUF_X1 U3 ( .A(n2), .Z(n11) );
  BUF_X1 U4 ( .A(n1), .Z(n8) );
  BUF_X1 U5 ( .A(n1), .Z(n7) );
  BUF_X1 U6 ( .A(n1), .Z(n6) );
  BUF_X1 U7 ( .A(n3), .Z(n14) );
  BUF_X1 U8 ( .A(n3), .Z(n13) );
  BUF_X1 U9 ( .A(n3), .Z(n12) );
  BUF_X1 U10 ( .A(n2), .Z(n10) );
  BUF_X1 U11 ( .A(n2), .Z(n9) );
  BUF_X1 U12 ( .A(sel), .Z(n3) );
  BUF_X1 U13 ( .A(sel), .Z(n2) );
  BUF_X1 U14 ( .A(sel), .Z(n1) );
  INV_X1 U15 ( .A(n53), .ZN(N4) );
  AOI22_X1 U16 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U17 ( .A(n54), .ZN(N5) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U19 ( .A(n55), .ZN(N6) );
  AOI22_X1 U20 ( .A1(port0[4]), .A2(n5), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U21 ( .A(n56), .ZN(N7) );
  AOI22_X1 U22 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U23 ( .A(n57), .ZN(N8) );
  AOI22_X1 U24 ( .A1(port0[6]), .A2(n5), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U25 ( .A(n58), .ZN(N9) );
  AOI22_X1 U26 ( .A1(port0[7]), .A2(n5), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U27 ( .A(n25), .ZN(N2) );
  AOI22_X1 U28 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  INV_X1 U29 ( .A(n48), .ZN(N3) );
  AOI22_X1 U30 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  INV_X1 U31 ( .A(n15), .ZN(N10) );
  AOI22_X1 U32 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U33 ( .A(n16), .ZN(N11) );
  AOI22_X1 U34 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U35 ( .A(n17), .ZN(N12) );
  AOI22_X1 U36 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U37 ( .A(n18), .ZN(N13) );
  AOI22_X1 U38 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U39 ( .A(n19), .ZN(N14) );
  AOI22_X1 U40 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U41 ( .A(n20), .ZN(N15) );
  AOI22_X1 U42 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U43 ( .A(n21), .ZN(N16) );
  AOI22_X1 U44 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U45 ( .A(n22), .ZN(N17) );
  AOI22_X1 U46 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  INV_X1 U47 ( .A(n23), .ZN(N18) );
  AOI22_X1 U48 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  INV_X1 U49 ( .A(n24), .ZN(N19) );
  AOI22_X1 U50 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U51 ( .A(n26), .ZN(N20) );
  AOI22_X1 U52 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  INV_X1 U53 ( .A(n51), .ZN(N32) );
  AOI22_X1 U54 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n7), .ZN(n51) );
  INV_X1 U55 ( .A(n27), .ZN(N21) );
  AOI22_X1 U56 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  INV_X1 U57 ( .A(n28), .ZN(N22) );
  AOI22_X1 U58 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U59 ( .A(n29), .ZN(N23) );
  AOI22_X1 U60 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  INV_X1 U61 ( .A(n30), .ZN(N24) );
  AOI22_X1 U62 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  INV_X1 U63 ( .A(n31), .ZN(N25) );
  AOI22_X1 U64 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  INV_X1 U65 ( .A(n32), .ZN(N26) );
  AOI22_X1 U66 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U67 ( .A(n33), .ZN(N27) );
  AOI22_X1 U68 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  INV_X1 U69 ( .A(n35), .ZN(N28) );
  AOI22_X1 U70 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  INV_X1 U71 ( .A(n47), .ZN(N29) );
  AOI22_X1 U72 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  INV_X1 U73 ( .A(n49), .ZN(N30) );
  AOI22_X1 U74 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U75 ( .A(n50), .ZN(N31) );
  AOI22_X1 U76 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  INV_X1 U77 ( .A(n52), .ZN(N33) );
  AOI22_X1 U78 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n7), .ZN(n52) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_15 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n5) );
  INV_X1 U2 ( .A(n14), .ZN(n4) );
  INV_X1 U3 ( .A(n57), .ZN(N8) );
  AOI22_X1 U4 ( .A1(port0[6]), .A2(n5), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U5 ( .A(n53), .ZN(N4) );
  AOI22_X1 U6 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U7 ( .A(n55), .ZN(N6) );
  AOI22_X1 U8 ( .A1(port0[4]), .A2(n5), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U9 ( .A(n56), .ZN(N7) );
  AOI22_X1 U10 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U11 ( .A(n54), .ZN(N5) );
  AOI22_X1 U12 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U13 ( .A(n58), .ZN(N9) );
  AOI22_X1 U14 ( .A1(port0[7]), .A2(n5), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U15 ( .A(n16), .ZN(N11) );
  AOI22_X1 U16 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U17 ( .A(n24), .ZN(N19) );
  AOI22_X1 U18 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U19 ( .A(n23), .ZN(N18) );
  AOI22_X1 U20 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  INV_X1 U21 ( .A(n25), .ZN(N2) );
  AOI22_X1 U22 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  INV_X1 U23 ( .A(n20), .ZN(N15) );
  AOI22_X1 U24 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U25 ( .A(n33), .ZN(N27) );
  AOI22_X1 U26 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  INV_X1 U27 ( .A(n19), .ZN(N14) );
  AOI22_X1 U28 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U29 ( .A(n17), .ZN(N12) );
  AOI22_X1 U30 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U31 ( .A(n28), .ZN(N22) );
  AOI22_X1 U32 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U33 ( .A(n29), .ZN(N23) );
  AOI22_X1 U34 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  INV_X1 U35 ( .A(n30), .ZN(N24) );
  AOI22_X1 U36 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  INV_X1 U37 ( .A(n26), .ZN(N20) );
  AOI22_X1 U38 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  INV_X1 U39 ( .A(n48), .ZN(N3) );
  AOI22_X1 U40 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  INV_X1 U41 ( .A(n21), .ZN(N16) );
  AOI22_X1 U42 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U43 ( .A(n49), .ZN(N30) );
  AOI22_X1 U44 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U45 ( .A(n50), .ZN(N31) );
  AOI22_X1 U46 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  INV_X1 U47 ( .A(n32), .ZN(N26) );
  AOI22_X1 U48 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U49 ( .A(n35), .ZN(N28) );
  AOI22_X1 U50 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  INV_X1 U51 ( .A(n15), .ZN(N10) );
  AOI22_X1 U52 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U53 ( .A(n18), .ZN(N13) );
  AOI22_X1 U54 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U55 ( .A(n22), .ZN(N17) );
  AOI22_X1 U56 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  INV_X1 U57 ( .A(n27), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  INV_X1 U59 ( .A(n31), .ZN(N25) );
  AOI22_X1 U60 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  INV_X1 U61 ( .A(n47), .ZN(N29) );
  AOI22_X1 U62 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  INV_X1 U63 ( .A(n51), .ZN(N32) );
  AOI22_X1 U64 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n7), .ZN(n51) );
  INV_X1 U65 ( .A(n52), .ZN(N33) );
  AOI22_X1 U66 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n7), .ZN(n52) );
  BUF_X1 U67 ( .A(n2), .Z(n11) );
  BUF_X1 U68 ( .A(n1), .Z(n8) );
  BUF_X1 U69 ( .A(n3), .Z(n12) );
  BUF_X1 U70 ( .A(n1), .Z(n6) );
  BUF_X1 U71 ( .A(n1), .Z(n7) );
  BUF_X1 U72 ( .A(n2), .Z(n10) );
  BUF_X1 U73 ( .A(n3), .Z(n14) );
  BUF_X1 U74 ( .A(n3), .Z(n13) );
  BUF_X1 U75 ( .A(n2), .Z(n9) );
  BUF_X1 U76 ( .A(sel), .Z(n2) );
  BUF_X1 U77 ( .A(sel), .Z(n3) );
  BUF_X1 U78 ( .A(sel), .Z(n1) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_14 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  AOI22_X1 U1 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n7), .ZN(n51) );
  AOI22_X1 U2 ( .A1(port0[7]), .A2(n5), .B1(n13), .B2(port1[7]), .ZN(n58) );
  AOI22_X1 U3 ( .A1(port0[31]), .A2(n4), .B1(port1[31]), .B2(n7), .ZN(n52) );
  AOI22_X1 U4 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17) );
  AOI22_X1 U5 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18) );
  AOI22_X1 U6 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  AOI22_X1 U7 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  AOI22_X1 U8 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26) );
  AOI22_X1 U9 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27) );
  AOI22_X1 U10 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  AOI22_X1 U11 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  AOI22_X1 U12 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  AOI22_X1 U13 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  AOI22_X1 U14 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n6), .ZN(n54) );
  AOI22_X1 U15 ( .A1(port0[6]), .A2(n5), .B1(port1[6]), .B2(n6), .ZN(n57) );
  AOI22_X1 U16 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U17 ( .A(n14), .ZN(n5) );
  INV_X1 U18 ( .A(n14), .ZN(n4) );
  AOI22_X1 U19 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  AOI22_X1 U20 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  AOI22_X1 U21 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  AOI22_X1 U22 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  AOI22_X1 U23 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  AOI22_X1 U24 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  AOI22_X1 U25 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n6), .ZN(n56) );
  AOI22_X1 U26 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  BUF_X1 U27 ( .A(n3), .Z(n14) );
  BUF_X1 U28 ( .A(n3), .Z(n12) );
  BUF_X1 U29 ( .A(n2), .Z(n11) );
  BUF_X1 U30 ( .A(n2), .Z(n10) );
  BUF_X1 U31 ( .A(n1), .Z(n7) );
  BUF_X1 U32 ( .A(n2), .Z(n9) );
  BUF_X1 U33 ( .A(n1), .Z(n8) );
  BUF_X1 U34 ( .A(n1), .Z(n6) );
  BUF_X1 U35 ( .A(n3), .Z(n13) );
  INV_X1 U36 ( .A(n25), .ZN(N2) );
  AOI22_X1 U37 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  AOI22_X1 U38 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  AOI22_X1 U39 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  AOI22_X1 U40 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  AOI22_X1 U41 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  AOI22_X1 U42 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U43 ( .A(n19), .ZN(N14) );
  INV_X1 U44 ( .A(n28), .ZN(N22) );
  INV_X1 U45 ( .A(n27), .ZN(N21) );
  INV_X1 U46 ( .A(n21), .ZN(N16) );
  INV_X1 U47 ( .A(n23), .ZN(N18) );
  INV_X1 U48 ( .A(n49), .ZN(N30) );
  INV_X1 U49 ( .A(n52), .ZN(N33) );
  INV_X1 U50 ( .A(n51), .ZN(N32) );
  INV_X1 U51 ( .A(n30), .ZN(N24) );
  INV_X1 U52 ( .A(n35), .ZN(N28) );
  INV_X1 U53 ( .A(n15), .ZN(N10) );
  INV_X1 U54 ( .A(n54), .ZN(N5) );
  INV_X1 U55 ( .A(n58), .ZN(N9) );
  INV_X1 U56 ( .A(n20), .ZN(N15) );
  INV_X1 U57 ( .A(n24), .ZN(N19) );
  INV_X1 U58 ( .A(n29), .ZN(N23) );
  INV_X1 U59 ( .A(n50), .ZN(N31) );
  INV_X1 U60 ( .A(n22), .ZN(N17) );
  INV_X1 U61 ( .A(n31), .ZN(N25) );
  INV_X1 U62 ( .A(n47), .ZN(N29) );
  INV_X1 U63 ( .A(n16), .ZN(N11) );
  INV_X1 U64 ( .A(n17), .ZN(N12) );
  INV_X1 U65 ( .A(n32), .ZN(N26) );
  INV_X1 U66 ( .A(n26), .ZN(N20) );
  INV_X1 U67 ( .A(n33), .ZN(N27) );
  INV_X1 U68 ( .A(n18), .ZN(N13) );
  AOI22_X1 U69 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U70 ( .A(n55), .ZN(N6) );
  INV_X1 U71 ( .A(n56), .ZN(N7) );
  INV_X1 U72 ( .A(n53), .ZN(N4) );
  INV_X1 U73 ( .A(n57), .ZN(N8) );
  INV_X1 U74 ( .A(n48), .ZN(N3) );
  AOI22_X1 U75 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  CLKBUF_X1 U76 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U77 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U78 ( .A(sel), .Z(n1) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_13 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n5) );
  INV_X1 U2 ( .A(n14), .ZN(n4) );
  BUF_X1 U3 ( .A(n1), .Z(n7) );
  BUF_X1 U4 ( .A(n3), .Z(n14) );
  BUF_X1 U5 ( .A(n3), .Z(n12) );
  BUF_X1 U6 ( .A(n2), .Z(n10) );
  BUF_X1 U7 ( .A(n2), .Z(n9) );
  BUF_X1 U8 ( .A(n1), .Z(n8) );
  BUF_X1 U9 ( .A(n1), .Z(n6) );
  BUF_X1 U10 ( .A(n3), .Z(n13) );
  BUF_X1 U11 ( .A(n2), .Z(n11) );
  INV_X1 U12 ( .A(n19), .ZN(N14) );
  INV_X1 U13 ( .A(n28), .ZN(N22) );
  INV_X1 U14 ( .A(n27), .ZN(N21) );
  INV_X1 U15 ( .A(n21), .ZN(N16) );
  INV_X1 U16 ( .A(n23), .ZN(N18) );
  INV_X1 U17 ( .A(n49), .ZN(N30) );
  INV_X1 U18 ( .A(n52), .ZN(N33) );
  INV_X1 U19 ( .A(n51), .ZN(N32) );
  INV_X1 U20 ( .A(n30), .ZN(N24) );
  INV_X1 U21 ( .A(n35), .ZN(N28) );
  INV_X1 U22 ( .A(n15), .ZN(N10) );
  INV_X1 U23 ( .A(n54), .ZN(N5) );
  INV_X1 U24 ( .A(n58), .ZN(N9) );
  INV_X1 U25 ( .A(n20), .ZN(N15) );
  INV_X1 U26 ( .A(n24), .ZN(N19) );
  INV_X1 U27 ( .A(n29), .ZN(N23) );
  INV_X1 U28 ( .A(n50), .ZN(N31) );
  INV_X1 U29 ( .A(n22), .ZN(N17) );
  INV_X1 U30 ( .A(n31), .ZN(N25) );
  INV_X1 U31 ( .A(n47), .ZN(N29) );
  INV_X1 U32 ( .A(n16), .ZN(N11) );
  INV_X1 U33 ( .A(n17), .ZN(N12) );
  INV_X1 U34 ( .A(n32), .ZN(N26) );
  INV_X1 U35 ( .A(n26), .ZN(N20) );
  INV_X1 U36 ( .A(n33), .ZN(N27) );
  INV_X1 U37 ( .A(n18), .ZN(N13) );
  INV_X1 U38 ( .A(n55), .ZN(N6) );
  INV_X1 U39 ( .A(n56), .ZN(N7) );
  INV_X1 U40 ( .A(n53), .ZN(N4) );
  INV_X1 U41 ( .A(n57), .ZN(N8) );
  INV_X1 U42 ( .A(n48), .ZN(N3) );
  CLKBUF_X1 U43 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U44 ( .A(sel), .Z(n1) );
  CLKBUF_X1 U45 ( .A(sel), .Z(n2) );
  AOI22_X1 U46 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  AOI22_X1 U47 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n6), .ZN(n55) );
  AOI22_X1 U48 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n6), .ZN(n56) );
  AOI22_X1 U49 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n7), .ZN(n51) );
  AOI22_X1 U50 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(n7), .ZN(n53) );
  AOI22_X1 U51 ( .A1(port0[7]), .A2(n5), .B1(n13), .B2(port1[7]), .ZN(n58) );
  AOI22_X1 U52 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n6), .ZN(n57) );
  AOI22_X1 U53 ( .A1(port0[31]), .A2(n4), .B1(port1[31]), .B2(n7), .ZN(n52) );
  AOI22_X1 U54 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  AOI22_X1 U55 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  AOI22_X1 U56 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  AOI22_X1 U57 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  AOI22_X1 U58 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  AOI22_X1 U59 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  AOI22_X1 U60 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  AOI22_X1 U61 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  AOI22_X1 U62 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  AOI22_X1 U63 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  AOI22_X1 U64 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  AOI22_X1 U65 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  AOI22_X1 U66 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  AOI22_X1 U67 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  AOI22_X1 U68 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  AOI22_X1 U69 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  AOI22_X1 U70 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  AOI22_X1 U71 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  AOI22_X1 U73 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  AOI22_X1 U75 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  AOI22_X1 U76 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  AOI22_X1 U77 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  INV_X1 U78 ( .A(n25), .ZN(N2) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_12 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n5) );
  INV_X1 U2 ( .A(n14), .ZN(n4) );
  BUF_X1 U3 ( .A(n3), .Z(n14) );
  BUF_X1 U4 ( .A(n3), .Z(n12) );
  BUF_X1 U5 ( .A(n2), .Z(n10) );
  BUF_X1 U6 ( .A(n1), .Z(n7) );
  BUF_X1 U7 ( .A(n2), .Z(n9) );
  BUF_X1 U8 ( .A(n1), .Z(n8) );
  BUF_X1 U9 ( .A(n1), .Z(n6) );
  BUF_X1 U10 ( .A(n3), .Z(n13) );
  BUF_X1 U11 ( .A(n2), .Z(n11) );
  CLKBUF_X1 U12 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U13 ( .A(sel), .Z(n2) );
  CLKBUF_X1 U14 ( .A(sel), .Z(n1) );
  INV_X1 U15 ( .A(n19), .ZN(N14) );
  AOI22_X1 U16 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U17 ( .A(n28), .ZN(N22) );
  AOI22_X1 U18 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U19 ( .A(n27), .ZN(N21) );
  AOI22_X1 U20 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  INV_X1 U21 ( .A(n21), .ZN(N16) );
  AOI22_X1 U22 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U23 ( .A(n23), .ZN(N18) );
  AOI22_X1 U24 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  INV_X1 U25 ( .A(n49), .ZN(N30) );
  AOI22_X1 U26 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U27 ( .A(n52), .ZN(N33) );
  AOI22_X1 U28 ( .A1(port0[31]), .A2(n4), .B1(port1[31]), .B2(n7), .ZN(n52) );
  INV_X1 U29 ( .A(n51), .ZN(N32) );
  AOI22_X1 U30 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n7), .ZN(n51) );
  INV_X1 U31 ( .A(n30), .ZN(N24) );
  AOI22_X1 U32 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  INV_X1 U33 ( .A(n35), .ZN(N28) );
  AOI22_X1 U34 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  INV_X1 U35 ( .A(n15), .ZN(N10) );
  AOI22_X1 U36 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U37 ( .A(n54), .ZN(N5) );
  AOI22_X1 U38 ( .A1(port0[3]), .A2(n4), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U39 ( .A(n58), .ZN(N9) );
  AOI22_X1 U40 ( .A1(port0[7]), .A2(n5), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U41 ( .A(n20), .ZN(N15) );
  AOI22_X1 U42 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U43 ( .A(n24), .ZN(N19) );
  AOI22_X1 U44 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U45 ( .A(n29), .ZN(N23) );
  AOI22_X1 U46 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  INV_X1 U47 ( .A(n50), .ZN(N31) );
  AOI22_X1 U48 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  INV_X1 U49 ( .A(n22), .ZN(N17) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  INV_X1 U51 ( .A(n31), .ZN(N25) );
  AOI22_X1 U52 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  INV_X1 U53 ( .A(n47), .ZN(N29) );
  AOI22_X1 U54 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  INV_X1 U55 ( .A(n16), .ZN(N11) );
  AOI22_X1 U56 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U57 ( .A(n17), .ZN(N12) );
  AOI22_X1 U58 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U59 ( .A(n32), .ZN(N26) );
  AOI22_X1 U60 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U61 ( .A(n26), .ZN(N20) );
  AOI22_X1 U62 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  INV_X1 U63 ( .A(n33), .ZN(N27) );
  AOI22_X1 U64 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  INV_X1 U65 ( .A(n18), .ZN(N13) );
  AOI22_X1 U66 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U67 ( .A(n55), .ZN(N6) );
  AOI22_X1 U68 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U69 ( .A(n56), .ZN(N7) );
  AOI22_X1 U70 ( .A1(port0[5]), .A2(n4), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U71 ( .A(n53), .ZN(N4) );
  AOI22_X1 U72 ( .A1(port0[2]), .A2(n5), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U73 ( .A(n57), .ZN(N8) );
  AOI22_X1 U74 ( .A1(port0[6]), .A2(n5), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U75 ( .A(n48), .ZN(N3) );
  AOI22_X1 U76 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  AOI22_X1 U77 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  INV_X1 U78 ( .A(n25), .ZN(N2) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_11 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  INV_X1 U3 ( .A(n53), .ZN(N4) );
  AOI22_X1 U4 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U5 ( .A(n54), .ZN(N5) );
  AOI22_X1 U6 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U7 ( .A(n55), .ZN(N6) );
  AOI22_X1 U8 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U9 ( .A(n56), .ZN(N7) );
  AOI22_X1 U10 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U11 ( .A(n57), .ZN(N8) );
  AOI22_X1 U12 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U13 ( .A(n51), .ZN(N32) );
  INV_X1 U14 ( .A(n52), .ZN(N33) );
  INV_X1 U15 ( .A(n58), .ZN(N9) );
  AOI22_X1 U16 ( .A1(port0[7]), .A2(n5), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U17 ( .A(n25), .ZN(N2) );
  AOI22_X1 U18 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  INV_X1 U19 ( .A(n48), .ZN(N3) );
  AOI22_X1 U20 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  INV_X1 U21 ( .A(n23), .ZN(N18) );
  INV_X1 U22 ( .A(n24), .ZN(N19) );
  INV_X1 U23 ( .A(n26), .ZN(N20) );
  INV_X1 U24 ( .A(n27), .ZN(N21) );
  INV_X1 U25 ( .A(n28), .ZN(N22) );
  INV_X1 U26 ( .A(n29), .ZN(N23) );
  INV_X1 U27 ( .A(n30), .ZN(N24) );
  INV_X1 U28 ( .A(n31), .ZN(N25) );
  INV_X1 U29 ( .A(n32), .ZN(N26) );
  INV_X1 U30 ( .A(n33), .ZN(N27) );
  INV_X1 U31 ( .A(n35), .ZN(N28) );
  INV_X1 U32 ( .A(n47), .ZN(N29) );
  INV_X1 U33 ( .A(n49), .ZN(N30) );
  INV_X1 U34 ( .A(n50), .ZN(N31) );
  BUF_X1 U35 ( .A(n1), .Z(n6) );
  BUF_X1 U36 ( .A(n3), .Z(n12) );
  BUF_X1 U37 ( .A(n2), .Z(n11) );
  BUF_X1 U38 ( .A(n2), .Z(n9) );
  BUF_X1 U39 ( .A(n1), .Z(n8) );
  BUF_X1 U40 ( .A(n2), .Z(n10) );
  BUF_X1 U41 ( .A(n1), .Z(n7) );
  BUF_X1 U42 ( .A(n3), .Z(n14) );
  BUF_X1 U43 ( .A(n3), .Z(n13) );
  INV_X1 U44 ( .A(n15), .ZN(N10) );
  AOI22_X1 U45 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U46 ( .A(n16), .ZN(N11) );
  AOI22_X1 U47 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U48 ( .A(n17), .ZN(N12) );
  AOI22_X1 U49 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U50 ( .A(n18), .ZN(N13) );
  AOI22_X1 U51 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U52 ( .A(n19), .ZN(N14) );
  AOI22_X1 U53 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U54 ( .A(n20), .ZN(N15) );
  AOI22_X1 U55 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U56 ( .A(n21), .ZN(N16) );
  AOI22_X1 U57 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U58 ( .A(n22), .ZN(N17) );
  AOI22_X1 U59 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  AOI22_X1 U60 ( .A1(port0[30]), .A2(n4), .B1(port1[30]), .B2(n7), .ZN(n51) );
  AOI22_X1 U61 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n7), .ZN(n52) );
  AOI22_X1 U62 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  AOI22_X1 U63 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  AOI22_X1 U64 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  AOI22_X1 U65 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  AOI22_X1 U66 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  AOI22_X1 U67 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  AOI22_X1 U68 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  AOI22_X1 U69 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  AOI22_X1 U70 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  AOI22_X1 U71 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  AOI22_X1 U73 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  AOI22_X1 U74 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  AOI22_X1 U75 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  BUF_X1 U76 ( .A(sel), .Z(n3) );
  BUF_X1 U77 ( .A(sel), .Z(n2) );
  BUF_X1 U78 ( .A(sel), .Z(n1) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_10 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  INV_X1 U3 ( .A(n53), .ZN(N4) );
  AOI22_X1 U4 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n7), .ZN(n53) );
  INV_X1 U5 ( .A(n54), .ZN(N5) );
  AOI22_X1 U6 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n54) );
  INV_X1 U7 ( .A(n55), .ZN(N6) );
  AOI22_X1 U8 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n6), .ZN(n55) );
  INV_X1 U9 ( .A(n56), .ZN(N7) );
  AOI22_X1 U10 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n56) );
  INV_X1 U11 ( .A(n57), .ZN(N8) );
  AOI22_X1 U12 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n6), .ZN(n57) );
  INV_X1 U13 ( .A(n51), .ZN(N32) );
  AOI22_X1 U14 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n7), .ZN(n51) );
  INV_X1 U15 ( .A(n52), .ZN(N33) );
  AOI22_X1 U16 ( .A1(port0[31]), .A2(n4), .B1(port1[31]), .B2(n7), .ZN(n52) );
  INV_X1 U17 ( .A(n58), .ZN(N9) );
  AOI22_X1 U18 ( .A1(port0[7]), .A2(n5), .B1(n13), .B2(port1[7]), .ZN(n58) );
  INV_X1 U19 ( .A(n25), .ZN(N2) );
  AOI22_X1 U20 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n25) );
  INV_X1 U21 ( .A(n48), .ZN(N3) );
  AOI22_X1 U22 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n48) );
  INV_X1 U23 ( .A(n23), .ZN(N18) );
  AOI22_X1 U24 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n23)
         );
  INV_X1 U25 ( .A(n24), .ZN(N19) );
  AOI22_X1 U26 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n24)
         );
  INV_X1 U27 ( .A(n26), .ZN(N20) );
  AOI22_X1 U28 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n26)
         );
  INV_X1 U29 ( .A(n27), .ZN(N21) );
  AOI22_X1 U30 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n27)
         );
  INV_X1 U31 ( .A(n28), .ZN(N22) );
  AOI22_X1 U32 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n28)
         );
  INV_X1 U33 ( .A(n29), .ZN(N23) );
  AOI22_X1 U34 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n29) );
  INV_X1 U35 ( .A(n30), .ZN(N24) );
  AOI22_X1 U36 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n30) );
  INV_X1 U37 ( .A(n31), .ZN(N25) );
  AOI22_X1 U38 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n31) );
  INV_X1 U39 ( .A(n32), .ZN(N26) );
  AOI22_X1 U40 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n32) );
  INV_X1 U41 ( .A(n33), .ZN(N27) );
  AOI22_X1 U42 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n33) );
  INV_X1 U43 ( .A(n35), .ZN(N28) );
  AOI22_X1 U44 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n35) );
  INV_X1 U45 ( .A(n47), .ZN(N29) );
  AOI22_X1 U46 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n47) );
  INV_X1 U47 ( .A(n49), .ZN(N30) );
  AOI22_X1 U48 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n49) );
  INV_X1 U49 ( .A(n50), .ZN(N31) );
  AOI22_X1 U50 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n50)
         );
  BUF_X1 U51 ( .A(n1), .Z(n6) );
  BUF_X1 U52 ( .A(n3), .Z(n12) );
  BUF_X1 U53 ( .A(n2), .Z(n11) );
  BUF_X1 U54 ( .A(n2), .Z(n9) );
  BUF_X1 U55 ( .A(n1), .Z(n8) );
  BUF_X1 U56 ( .A(n2), .Z(n10) );
  BUF_X1 U57 ( .A(n1), .Z(n7) );
  BUF_X1 U58 ( .A(n3), .Z(n14) );
  BUF_X1 U59 ( .A(n3), .Z(n13) );
  INV_X1 U60 ( .A(n15), .ZN(N10) );
  AOI22_X1 U61 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n15) );
  INV_X1 U62 ( .A(n16), .ZN(N11) );
  AOI22_X1 U63 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n16) );
  INV_X1 U64 ( .A(n17), .ZN(N12) );
  AOI22_X1 U65 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n17)
         );
  INV_X1 U66 ( .A(n18), .ZN(N13) );
  AOI22_X1 U67 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n18)
         );
  INV_X1 U68 ( .A(n19), .ZN(N14) );
  AOI22_X1 U69 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n19)
         );
  INV_X1 U70 ( .A(n20), .ZN(N15) );
  AOI22_X1 U71 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n20)
         );
  INV_X1 U72 ( .A(n21), .ZN(N16) );
  AOI22_X1 U73 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n21)
         );
  INV_X1 U74 ( .A(n22), .ZN(N17) );
  AOI22_X1 U75 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n22)
         );
  BUF_X1 U76 ( .A(sel), .Z(n3) );
  BUF_X1 U77 ( .A(sel), .Z(n2) );
  BUF_X1 U78 ( .A(sel), .Z(n1) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_9 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n57, n58, n59, net132973, net132971, net132967,
         net132965, net132963, net132961, net132959, net132957, net132955,
         net132953, net132979, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25,
         n26, n27, n28, n29, n30, n31, n32, n33;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  AOI22_X1 U1 ( .A1(port0[0]), .A2(net132953), .B1(port1[0]), .B2(n2), .ZN(n1)
         );
  INV_X1 U2 ( .A(n1), .ZN(N2) );
  BUF_X1 U3 ( .A(n4), .Z(n2) );
  AOI22_X1 U4 ( .A1(port0[15]), .A2(net132953), .B1(port1[15]), .B2(n2), .ZN(
        n59) );
  AOI22_X1 U5 ( .A1(port0[16]), .A2(net132953), .B1(port1[16]), .B2(n2), .ZN(
        n58) );
  AOI22_X1 U6 ( .A1(port0[17]), .A2(net132953), .B1(port1[17]), .B2(n2), .ZN(
        n57) );
  CLKBUF_X1 U7 ( .A(sel), .Z(n4) );
  BUF_X1 U8 ( .A(n4), .Z(net132967) );
  BUF_X1 U9 ( .A(n4), .Z(net132965) );
  INV_X1 U10 ( .A(n3), .ZN(net132953) );
  BUF_X1 U11 ( .A(n5), .Z(n3) );
  INV_X1 U12 ( .A(n3), .ZN(net132955) );
  INV_X1 U13 ( .A(n3), .ZN(net132957) );
  BUF_X1 U14 ( .A(sel), .Z(n5) );
  CLKBUF_X1 U15 ( .A(n5), .Z(net132971) );
  CLKBUF_X1 U16 ( .A(n5), .Z(net132973) );
  CLKBUF_X1 U17 ( .A(sel), .Z(net132979) );
  CLKBUF_X1 U18 ( .A(net132979), .Z(net132959) );
  INV_X1 U19 ( .A(n33), .ZN(N9) );
  INV_X1 U20 ( .A(n21), .ZN(N28) );
  INV_X1 U21 ( .A(n23), .ZN(N3) );
  AOI22_X1 U22 ( .A1(port0[1]), .A2(net132955), .B1(port1[1]), .B2(net132963), 
        .ZN(n23) );
  INV_X1 U23 ( .A(n17), .ZN(N24) );
  INV_X1 U24 ( .A(n16), .ZN(N23) );
  INV_X1 U25 ( .A(n25), .ZN(N31) );
  INV_X1 U26 ( .A(n22), .ZN(N29) );
  INV_X1 U27 ( .A(n24), .ZN(N30) );
  INV_X1 U28 ( .A(n20), .ZN(N27) );
  INV_X1 U29 ( .A(n18), .ZN(N25) );
  INV_X1 U30 ( .A(n14), .ZN(N21) );
  INV_X1 U31 ( .A(n15), .ZN(N22) );
  INV_X1 U32 ( .A(n30), .ZN(N6) );
  AOI22_X1 U33 ( .A1(port0[4]), .A2(net132957), .B1(port1[4]), .B2(net132959), 
        .ZN(n30) );
  INV_X1 U34 ( .A(n28), .ZN(N4) );
  AOI22_X1 U35 ( .A1(port0[2]), .A2(net132957), .B1(port1[2]), .B2(net132961), 
        .ZN(n28) );
  INV_X1 U36 ( .A(n29), .ZN(N5) );
  AOI22_X1 U37 ( .A1(port0[3]), .A2(net132957), .B1(port1[3]), .B2(net132959), 
        .ZN(n29) );
  INV_X1 U38 ( .A(n12), .ZN(N16) );
  INV_X1 U39 ( .A(n10), .ZN(N14) );
  AOI22_X1 U40 ( .A1(port0[12]), .A2(net132953), .B1(port1[12]), .B2(net132971), .ZN(n10) );
  INV_X1 U41 ( .A(n59), .ZN(N17) );
  INV_X1 U42 ( .A(n31), .ZN(N7) );
  AOI22_X1 U43 ( .A1(port0[5]), .A2(net132957), .B1(port1[5]), .B2(net132959), 
        .ZN(n31) );
  INV_X1 U44 ( .A(n13), .ZN(N20) );
  INV_X1 U45 ( .A(n6), .ZN(N10) );
  INV_X1 U46 ( .A(n7), .ZN(N11) );
  INV_X1 U47 ( .A(n9), .ZN(N13) );
  AOI22_X1 U48 ( .A1(port0[11]), .A2(net132953), .B1(port1[11]), .B2(net132971), .ZN(n9) );
  INV_X1 U49 ( .A(n11), .ZN(N15) );
  INV_X1 U50 ( .A(n57), .ZN(N19) );
  INV_X1 U51 ( .A(n58), .ZN(N18) );
  INV_X1 U52 ( .A(n8), .ZN(N12) );
  INV_X1 U53 ( .A(n32), .ZN(N8) );
  AOI22_X1 U54 ( .A1(port0[6]), .A2(net132957), .B1(port1[6]), .B2(net132959), 
        .ZN(n32) );
  BUF_X1 U55 ( .A(net132979), .Z(net132961) );
  CLKBUF_X1 U56 ( .A(net132979), .Z(net132963) );
  AOI22_X1 U57 ( .A1(port0[22]), .A2(net132955), .B1(port1[22]), .B2(net132965), .ZN(n17) );
  AOI22_X1 U58 ( .A1(port0[13]), .A2(net132953), .B1(port1[13]), .B2(net132971), .ZN(n11) );
  AOI22_X1 U59 ( .A1(port0[10]), .A2(net132953), .B1(port1[10]), .B2(net132973), .ZN(n8) );
  AOI22_X1 U60 ( .A1(port0[14]), .A2(net132953), .B1(port1[14]), .B2(net132971), .ZN(n12) );
  AOI22_X1 U61 ( .A1(port0[8]), .A2(net132953), .B1(port1[8]), .B2(net132973), 
        .ZN(n6) );
  INV_X1 U62 ( .A(n19), .ZN(N26) );
  AOI22_X1 U63 ( .A1(port0[21]), .A2(net132955), .B1(port1[21]), .B2(net132965), .ZN(n16) );
  AOI22_X1 U64 ( .A1(port0[20]), .A2(net132955), .B1(port1[20]), .B2(net132967), .ZN(n15) );
  AOI22_X1 U65 ( .A1(port0[23]), .A2(net132955), .B1(port1[23]), .B2(net132965), .ZN(n18) );
  AOI22_X1 U66 ( .A1(port0[9]), .A2(net132953), .B1(port1[9]), .B2(net132973), 
        .ZN(n7) );
  INV_X1 U67 ( .A(n26), .ZN(N32) );
  AOI22_X1 U68 ( .A1(port0[7]), .A2(net132957), .B1(net132973), .B2(port1[7]), 
        .ZN(n33) );
  AOI22_X1 U69 ( .A1(port0[29]), .A2(net132955), .B1(port1[29]), .B2(net132967), .ZN(n25) );
  AOI22_X1 U70 ( .A1(port0[28]), .A2(net132955), .B1(port1[28]), .B2(net132961), .ZN(n24) );
  AOI22_X1 U71 ( .A1(port0[18]), .A2(net132953), .B1(port1[18]), .B2(net132967), .ZN(n13) );
  AOI22_X1 U72 ( .A1(port0[19]), .A2(net132955), .B1(port1[19]), .B2(net132967), .ZN(n14) );
  AOI22_X1 U73 ( .A1(port0[30]), .A2(net132957), .B1(port1[30]), .B2(net132961), .ZN(n26) );
  AOI22_X1 U74 ( .A1(port0[26]), .A2(net132955), .B1(port1[26]), .B2(net132963), .ZN(n21) );
  AOI22_X1 U75 ( .A1(port0[27]), .A2(net132955), .B1(port1[27]), .B2(net132963), .ZN(n22) );
  AOI22_X1 U76 ( .A1(port0[25]), .A2(net132955), .B1(port1[25]), .B2(net132963), .ZN(n20) );
  AOI22_X1 U77 ( .A1(port0[24]), .A2(net132955), .B1(port1[24]), .B2(net132965), .ZN(n19) );
  INV_X1 U78 ( .A(n27), .ZN(N33) );
  AOI22_X1 U79 ( .A1(port0[31]), .A2(net132957), .B1(port1[31]), .B2(net132961), .ZN(n27) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_8 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, n57, n58, n59, net132943, net132941, net132937, net132935,
         net132933, net132931, net132929, net132927, net132925, net132923,
         net132947, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;

  MUX2_X2 U1 ( .A(port1[25]), .B(port0[25]), .S(net132927), .Z(N27) );
  MUX2_X2 U2 ( .A(port0[3]), .B(port1[3]), .S(sel), .Z(N5) );
  NAND2_X1 U3 ( .A1(port0[31]), .A2(net132927), .ZN(n1) );
  NAND2_X1 U4 ( .A1(port1[31]), .A2(net132931), .ZN(n2) );
  NAND2_X1 U5 ( .A1(n2), .A2(n1), .ZN(portY[31]) );
  MUX2_X1 U6 ( .A(port0[0]), .B(port1[0]), .S(sel), .Z(N2) );
  BUF_X1 U7 ( .A(n6), .Z(n4) );
  AOI22_X1 U8 ( .A1(port0[17]), .A2(net132923), .B1(port1[17]), .B2(n4), .ZN(
        n57) );
  AOI22_X1 U9 ( .A1(port0[16]), .A2(net132923), .B1(port1[16]), .B2(n4), .ZN(
        n58) );
  AOI22_X1 U10 ( .A1(port0[15]), .A2(net132923), .B1(port1[15]), .B2(n4), .ZN(
        n59) );
  CLKBUF_X1 U11 ( .A(sel), .Z(n6) );
  BUF_X1 U12 ( .A(n6), .Z(net132935) );
  BUF_X1 U13 ( .A(n6), .Z(net132937) );
  INV_X1 U14 ( .A(n5), .ZN(net132923) );
  BUF_X1 U15 ( .A(n7), .Z(n5) );
  INV_X1 U16 ( .A(n5), .ZN(net132925) );
  INV_X1 U17 ( .A(n5), .ZN(net132927) );
  BUF_X1 U18 ( .A(sel), .Z(n7) );
  CLKBUF_X1 U19 ( .A(n7), .Z(net132943) );
  BUF_X1 U20 ( .A(n7), .Z(net132941) );
  CLKBUF_X1 U21 ( .A(sel), .Z(net132947) );
  CLKBUF_X1 U22 ( .A(net132947), .Z(net132929) );
  CLKBUF_X1 U23 ( .A(net132947), .Z(net132933) );
  INV_X1 U24 ( .A(n32), .ZN(N9) );
  AOI22_X1 U25 ( .A1(port0[30]), .A2(net132927), .B1(port1[30]), .B2(net132931), .ZN(n27) );
  INV_X1 U26 ( .A(n22), .ZN(N28) );
  AOI22_X1 U27 ( .A1(port0[26]), .A2(net132925), .B1(port1[26]), .B2(net132933), .ZN(n22) );
  INV_X1 U28 ( .A(n24), .ZN(N3) );
  AOI22_X1 U29 ( .A1(port0[1]), .A2(net132925), .B1(port1[1]), .B2(net132933), 
        .ZN(n24) );
  INV_X1 U30 ( .A(n19), .ZN(N24) );
  AOI22_X1 U31 ( .A1(port0[22]), .A2(net132925), .B1(port1[22]), .B2(net132935), .ZN(n19) );
  INV_X1 U32 ( .A(n18), .ZN(N23) );
  AOI22_X1 U33 ( .A1(port0[21]), .A2(net132925), .B1(port1[21]), .B2(net132935), .ZN(n18) );
  INV_X1 U34 ( .A(n26), .ZN(N31) );
  AOI22_X1 U35 ( .A1(port0[29]), .A2(net132925), .B1(port1[29]), .B2(net132937), .ZN(n26) );
  INV_X1 U36 ( .A(n23), .ZN(N29) );
  AOI22_X1 U37 ( .A1(port0[27]), .A2(net132925), .B1(port1[27]), .B2(net132933), .ZN(n23) );
  INV_X1 U38 ( .A(n25), .ZN(N30) );
  AOI22_X1 U39 ( .A1(port0[28]), .A2(net132925), .B1(port1[28]), .B2(net132931), .ZN(n25) );
  INV_X1 U40 ( .A(n20), .ZN(N25) );
  AOI22_X1 U41 ( .A1(port0[23]), .A2(net132925), .B1(port1[23]), .B2(net132935), .ZN(n20) );
  INV_X1 U42 ( .A(n16), .ZN(N21) );
  AOI22_X1 U43 ( .A1(port0[19]), .A2(net132925), .B1(port1[19]), .B2(net132937), .ZN(n16) );
  INV_X1 U44 ( .A(n21), .ZN(N26) );
  AOI22_X1 U45 ( .A1(port0[24]), .A2(net132925), .B1(port1[24]), .B2(net132935), .ZN(n21) );
  INV_X1 U46 ( .A(n17), .ZN(N22) );
  AOI22_X1 U47 ( .A1(port0[20]), .A2(net132925), .B1(port1[20]), .B2(net132937), .ZN(n17) );
  INV_X1 U48 ( .A(n29), .ZN(N6) );
  AOI22_X1 U49 ( .A1(port0[4]), .A2(net132927), .B1(port1[4]), .B2(net132929), 
        .ZN(n29) );
  INV_X1 U50 ( .A(n28), .ZN(N4) );
  AOI22_X1 U51 ( .A1(port0[2]), .A2(net132927), .B1(port1[2]), .B2(net132931), 
        .ZN(n28) );
  INV_X1 U52 ( .A(n14), .ZN(N16) );
  AOI22_X1 U53 ( .A1(port0[14]), .A2(net132923), .B1(port1[14]), .B2(net132941), .ZN(n14) );
  INV_X1 U54 ( .A(n12), .ZN(N14) );
  AOI22_X1 U55 ( .A1(port0[12]), .A2(net132923), .B1(port1[12]), .B2(net132941), .ZN(n12) );
  INV_X1 U56 ( .A(n59), .ZN(N17) );
  INV_X1 U57 ( .A(n30), .ZN(N7) );
  AOI22_X1 U58 ( .A1(port0[5]), .A2(net132927), .B1(port1[5]), .B2(net132929), 
        .ZN(n30) );
  INV_X1 U59 ( .A(n15), .ZN(N20) );
  AOI22_X1 U60 ( .A1(port0[18]), .A2(net132923), .B1(port1[18]), .B2(net132937), .ZN(n15) );
  INV_X1 U61 ( .A(n8), .ZN(N10) );
  AOI22_X1 U62 ( .A1(port0[8]), .A2(net132923), .B1(port1[8]), .B2(net132943), 
        .ZN(n8) );
  INV_X1 U63 ( .A(n9), .ZN(N11) );
  AOI22_X1 U64 ( .A1(port0[9]), .A2(net132923), .B1(port1[9]), .B2(net132943), 
        .ZN(n9) );
  INV_X1 U65 ( .A(n11), .ZN(N13) );
  AOI22_X1 U66 ( .A1(port0[11]), .A2(net132923), .B1(port1[11]), .B2(net132941), .ZN(n11) );
  INV_X1 U67 ( .A(n13), .ZN(N15) );
  AOI22_X1 U68 ( .A1(port0[13]), .A2(net132923), .B1(port1[13]), .B2(net132941), .ZN(n13) );
  INV_X1 U69 ( .A(n57), .ZN(N19) );
  INV_X1 U70 ( .A(n58), .ZN(N18) );
  INV_X1 U71 ( .A(n10), .ZN(N12) );
  AOI22_X1 U72 ( .A1(port0[10]), .A2(net132923), .B1(port1[10]), .B2(net132943), .ZN(n10) );
  INV_X1 U73 ( .A(n31), .ZN(N8) );
  AOI22_X1 U74 ( .A1(port0[6]), .A2(net132927), .B1(port1[6]), .B2(net132929), 
        .ZN(n31) );
  BUF_X1 U75 ( .A(net132947), .Z(net132931) );
  INV_X1 U76 ( .A(n27), .ZN(N32) );
  AOI22_X1 U77 ( .A1(port0[7]), .A2(net132927), .B1(net132943), .B2(port1[7]), 
        .ZN(n32) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_3 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n38, n39, n40;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  BUF_X4 U1 ( .A(sel), .Z(n5) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n4) );
  INV_X2 U3 ( .A(sel), .ZN(n3) );
  INV_X1 U4 ( .A(n26), .ZN(N29) );
  INV_X1 U5 ( .A(n25), .ZN(N28) );
  INV_X1 U6 ( .A(n24), .ZN(N27) );
  AOI22_X1 U7 ( .A1(port0[26]), .A2(n3), .B1(port1[26]), .B2(n5), .ZN(n25) );
  AOI22_X1 U8 ( .A1(port0[28]), .A2(n3), .B1(port1[28]), .B2(n5), .ZN(n28) );
  AOI22_X1 U9 ( .A1(port0[27]), .A2(n3), .B1(port1[27]), .B2(n5), .ZN(n26) );
  AOI22_X1 U10 ( .A1(port0[29]), .A2(n3), .B1(port1[29]), .B2(n4), .ZN(n29) );
  AOI22_X1 U11 ( .A1(port0[25]), .A2(n3), .B1(port1[25]), .B2(n5), .ZN(n24) );
  INV_X1 U12 ( .A(n29), .ZN(N31) );
  INV_X1 U13 ( .A(n28), .ZN(N30) );
  INV_X1 U14 ( .A(n17), .ZN(N20) );
  INV_X1 U15 ( .A(n23), .ZN(N26) );
  INV_X1 U16 ( .A(n13), .ZN(N17) );
  INV_X1 U17 ( .A(n14), .ZN(N18) );
  INV_X1 U18 ( .A(n19), .ZN(N22) );
  INV_X1 U19 ( .A(n15), .ZN(N19) );
  INV_X1 U20 ( .A(n12), .ZN(N16) );
  INV_X1 U21 ( .A(n18), .ZN(N21) );
  INV_X1 U22 ( .A(n11), .ZN(N15) );
  INV_X1 U23 ( .A(n8), .ZN(N12) );
  INV_X1 U24 ( .A(n21), .ZN(N24) );
  INV_X1 U25 ( .A(n5), .ZN(n2) );
  INV_X1 U26 ( .A(n22), .ZN(N25) );
  AOI22_X1 U27 ( .A1(port0[24]), .A2(n3), .B1(port1[24]), .B2(n5), .ZN(n23) );
  AOI22_X1 U28 ( .A1(port0[23]), .A2(n3), .B1(port1[23]), .B2(n4), .ZN(n22) );
  AOI22_X1 U29 ( .A1(port0[21]), .A2(n3), .B1(port1[21]), .B2(n4), .ZN(n20) );
  AOI22_X1 U30 ( .A1(port0[22]), .A2(n3), .B1(port1[22]), .B2(n5), .ZN(n21) );
  INV_X1 U31 ( .A(n20), .ZN(N23) );
  INV_X1 U32 ( .A(n10), .ZN(N14) );
  INV_X1 U33 ( .A(n9), .ZN(N13) );
  INV_X1 U34 ( .A(n7), .ZN(N11) );
  INV_X1 U35 ( .A(n33), .ZN(N5) );
  INV_X1 U36 ( .A(n39), .ZN(N8) );
  INV_X1 U37 ( .A(n27), .ZN(N3) );
  INV_X1 U38 ( .A(n16), .ZN(N2) );
  INV_X1 U39 ( .A(n6), .ZN(N10) );
  INV_X1 U40 ( .A(n38), .ZN(N7) );
  INV_X1 U41 ( .A(n35), .ZN(N6) );
  INV_X1 U42 ( .A(n32), .ZN(N4) );
  INV_X1 U43 ( .A(n40), .ZN(N9) );
  AOI22_X1 U44 ( .A1(port0[16]), .A2(n2), .B1(port1[16]), .B2(n5), .ZN(n14) );
  AOI22_X1 U45 ( .A1(port0[20]), .A2(n3), .B1(port1[20]), .B2(n4), .ZN(n19) );
  AOI22_X1 U46 ( .A1(port0[15]), .A2(n2), .B1(port1[15]), .B2(n5), .ZN(n13) );
  AOI22_X1 U47 ( .A1(port0[18]), .A2(n2), .B1(port1[18]), .B2(n4), .ZN(n17) );
  AOI22_X1 U48 ( .A1(port0[17]), .A2(n2), .B1(port1[17]), .B2(n5), .ZN(n15) );
  AOI22_X1 U49 ( .A1(port0[19]), .A2(n3), .B1(port1[19]), .B2(n4), .ZN(n18) );
  AOI22_X1 U50 ( .A1(port0[13]), .A2(n2), .B1(port1[13]), .B2(n5), .ZN(n11) );
  AOI22_X1 U51 ( .A1(port0[12]), .A2(n2), .B1(port1[12]), .B2(n5), .ZN(n10) );
  AOI22_X1 U52 ( .A1(port0[10]), .A2(n2), .B1(port1[10]), .B2(n5), .ZN(n8) );
  AOI22_X1 U53 ( .A1(port0[14]), .A2(n2), .B1(port1[14]), .B2(n5), .ZN(n12) );
  AOI22_X1 U54 ( .A1(port0[11]), .A2(n2), .B1(port1[11]), .B2(n5), .ZN(n9) );
  AOI22_X1 U55 ( .A1(port0[9]), .A2(n2), .B1(port1[9]), .B2(n5), .ZN(n7) );
  AOI22_X1 U56 ( .A1(port0[6]), .A2(n2), .B1(port1[6]), .B2(n5), .ZN(n39) );
  AOI22_X1 U57 ( .A1(port0[2]), .A2(n2), .B1(port1[2]), .B2(n5), .ZN(n32) );
  AOI22_X1 U58 ( .A1(port0[4]), .A2(n2), .B1(port1[4]), .B2(n5), .ZN(n35) );
  AOI22_X1 U59 ( .A1(port0[5]), .A2(n2), .B1(port1[5]), .B2(n5), .ZN(n38) );
  AOI22_X1 U60 ( .A1(port0[3]), .A2(n2), .B1(port1[3]), .B2(n5), .ZN(n33) );
  AOI22_X1 U61 ( .A1(port0[7]), .A2(n2), .B1(n5), .B2(port1[7]), .ZN(n40) );
  AOI22_X1 U62 ( .A1(port0[0]), .A2(n2), .B1(port1[0]), .B2(n5), .ZN(n16) );
  AOI22_X1 U63 ( .A1(port0[1]), .A2(n3), .B1(port1[1]), .B2(n5), .ZN(n27) );
  AOI22_X1 U64 ( .A1(port0[8]), .A2(n2), .B1(port1[8]), .B2(n5), .ZN(n6) );
  CLKBUF_X1 U65 ( .A(sel), .Z(n1) );
  AOI22_X1 U66 ( .A1(port0[30]), .A2(n3), .B1(port1[30]), .B2(n1), .ZN(n30) );
  AOI22_X1 U67 ( .A1(port0[31]), .A2(n3), .B1(port1[31]), .B2(n1), .ZN(n31) );
  INV_X1 U68 ( .A(n30), .ZN(N32) );
  INV_X1 U69 ( .A(n31), .ZN(N33) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_2 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13,
         n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27,
         n28, n29, n30, n31, n32, n33, n35, n40, n41, n42, n43, n44;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  BUF_X1 U1 ( .A(sel), .Z(n2) );
  BUF_X2 U2 ( .A(n2), .Z(n6) );
  BUF_X2 U3 ( .A(n1), .Z(n5) );
  INV_X2 U4 ( .A(n2), .ZN(n4) );
  INV_X1 U5 ( .A(n28), .ZN(N29) );
  INV_X1 U6 ( .A(n27), .ZN(N28) );
  INV_X1 U7 ( .A(n26), .ZN(N27) );
  AOI22_X1 U8 ( .A1(port0[26]), .A2(n4), .B1(port1[26]), .B2(n7), .ZN(n27) );
  AOI22_X1 U9 ( .A1(port0[28]), .A2(n4), .B1(port1[28]), .B2(n6), .ZN(n30) );
  AOI22_X1 U10 ( .A1(port0[25]), .A2(n4), .B1(port1[25]), .B2(n7), .ZN(n26) );
  AOI22_X1 U11 ( .A1(port0[29]), .A2(n4), .B1(port1[29]), .B2(n6), .ZN(n31) );
  AOI22_X1 U12 ( .A1(port0[27]), .A2(n4), .B1(port1[27]), .B2(n5), .ZN(n28) );
  INV_X1 U13 ( .A(n31), .ZN(N31) );
  INV_X1 U14 ( .A(n30), .ZN(N30) );
  INV_X1 U15 ( .A(n19), .ZN(N20) );
  INV_X1 U16 ( .A(n25), .ZN(N26) );
  INV_X1 U17 ( .A(n15), .ZN(N17) );
  INV_X1 U18 ( .A(n16), .ZN(N18) );
  INV_X1 U19 ( .A(n21), .ZN(N22) );
  INV_X1 U20 ( .A(n17), .ZN(N19) );
  INV_X1 U21 ( .A(n14), .ZN(N16) );
  INV_X1 U22 ( .A(n20), .ZN(N21) );
  INV_X1 U23 ( .A(n13), .ZN(N15) );
  INV_X1 U24 ( .A(n10), .ZN(N12) );
  INV_X1 U25 ( .A(n23), .ZN(N24) );
  INV_X1 U26 ( .A(n5), .ZN(n3) );
  INV_X1 U27 ( .A(n24), .ZN(N25) );
  INV_X1 U28 ( .A(n22), .ZN(N23) );
  INV_X1 U29 ( .A(n12), .ZN(N14) );
  INV_X1 U30 ( .A(n11), .ZN(N13) );
  INV_X1 U31 ( .A(n9), .ZN(N11) );
  INV_X1 U32 ( .A(n40), .ZN(N5) );
  INV_X1 U33 ( .A(n43), .ZN(N8) );
  INV_X1 U34 ( .A(n29), .ZN(N3) );
  INV_X1 U35 ( .A(n18), .ZN(N2) );
  INV_X1 U36 ( .A(n8), .ZN(N10) );
  INV_X1 U37 ( .A(n42), .ZN(N7) );
  INV_X1 U38 ( .A(n41), .ZN(N6) );
  INV_X1 U39 ( .A(n35), .ZN(N4) );
  INV_X1 U40 ( .A(n44), .ZN(N9) );
  AOI22_X1 U41 ( .A1(port0[16]), .A2(n3), .B1(port1[16]), .B2(n7), .ZN(n16) );
  AOI22_X1 U42 ( .A1(port0[20]), .A2(n4), .B1(port1[20]), .B2(n5), .ZN(n21) );
  AOI22_X1 U43 ( .A1(port0[15]), .A2(n3), .B1(port1[15]), .B2(n7), .ZN(n15) );
  AOI22_X1 U44 ( .A1(port0[18]), .A2(n3), .B1(port1[18]), .B2(n7), .ZN(n19) );
  AOI22_X1 U45 ( .A1(port0[17]), .A2(n3), .B1(port1[17]), .B2(n7), .ZN(n17) );
  AOI22_X1 U46 ( .A1(port0[19]), .A2(n4), .B1(port1[19]), .B2(n7), .ZN(n20) );
  AOI22_X1 U47 ( .A1(port0[10]), .A2(n3), .B1(port1[10]), .B2(n7), .ZN(n10) );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n3), .B1(port1[14]), .B2(n7), .ZN(n14) );
  AOI22_X1 U49 ( .A1(port0[11]), .A2(n3), .B1(port1[11]), .B2(n7), .ZN(n11) );
  CLKBUF_X1 U50 ( .A(n2), .Z(n7) );
  AOI22_X1 U51 ( .A1(port0[13]), .A2(n3), .B1(port1[13]), .B2(n7), .ZN(n13) );
  AOI22_X1 U52 ( .A1(port0[23]), .A2(n4), .B1(port1[23]), .B2(n6), .ZN(n24) );
  AOI22_X1 U53 ( .A1(port0[21]), .A2(n4), .B1(port1[21]), .B2(n6), .ZN(n22) );
  AOI22_X1 U54 ( .A1(port0[22]), .A2(n4), .B1(port1[22]), .B2(n6), .ZN(n23) );
  AOI22_X1 U55 ( .A1(port0[24]), .A2(n4), .B1(port1[24]), .B2(n6), .ZN(n25) );
  AOI22_X1 U56 ( .A1(port0[12]), .A2(n3), .B1(port1[12]), .B2(n7), .ZN(n12) );
  AOI22_X1 U57 ( .A1(port0[9]), .A2(n3), .B1(port1[9]), .B2(n7), .ZN(n9) );
  AOI22_X1 U58 ( .A1(port0[2]), .A2(n3), .B1(port1[2]), .B2(n7), .ZN(n35) );
  AOI22_X1 U59 ( .A1(port0[4]), .A2(n3), .B1(port1[4]), .B2(n5), .ZN(n41) );
  AOI22_X1 U60 ( .A1(port0[5]), .A2(n3), .B1(port1[5]), .B2(n5), .ZN(n42) );
  AOI22_X1 U61 ( .A1(port0[3]), .A2(n3), .B1(port1[3]), .B2(n5), .ZN(n40) );
  AOI22_X1 U62 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n7), .ZN(n29) );
  AOI22_X1 U63 ( .A1(port0[7]), .A2(n3), .B1(n7), .B2(port1[7]), .ZN(n44) );
  AOI22_X1 U64 ( .A1(port0[8]), .A2(n3), .B1(port1[8]), .B2(n7), .ZN(n8) );
  AOI22_X1 U65 ( .A1(port0[6]), .A2(n3), .B1(port1[6]), .B2(n5), .ZN(n43) );
  AOI22_X1 U66 ( .A1(port0[0]), .A2(n3), .B1(port1[0]), .B2(n7), .ZN(n18) );
  CLKBUF_X1 U67 ( .A(sel), .Z(n1) );
  AOI22_X1 U68 ( .A1(port0[31]), .A2(n4), .B1(port1[31]), .B2(n1), .ZN(n33) );
  INV_X1 U69 ( .A(n32), .ZN(N32) );
  INV_X1 U70 ( .A(n33), .ZN(N33) );
  AOI22_X1 U71 ( .A1(port0[30]), .A2(n4), .B1(port1[30]), .B2(n1), .ZN(n32) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_1 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N33, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n35, n42, n44, n45, n46, n47, n48, n49, n50,
         n51;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[31] = N33;

  INV_X2 U31 ( .A(n29), .ZN(N25) );
  BUF_X2 U1 ( .A(n5), .Z(n12) );
  INV_X4 U2 ( .A(n12), .ZN(n6) );
  INV_X1 U3 ( .A(n26), .ZN(N22) );
  INV_X1 U4 ( .A(n42), .ZN(N30) );
  INV_X1 U5 ( .A(n22), .ZN(N19) );
  INV_X1 U6 ( .A(n27), .ZN(N23) );
  BUF_X1 U7 ( .A(n4), .Z(n7) );
  INV_X1 U8 ( .A(n24), .ZN(N20) );
  INV_X1 U9 ( .A(n28), .ZN(N24) );
  INV_X1 U10 ( .A(n32), .ZN(N28) );
  INV_X1 U11 ( .A(n25), .ZN(N21) );
  NAND2_X1 U12 ( .A1(n2), .A2(n3), .ZN(portY[30]) );
  NAND2_X1 U13 ( .A1(port0[30]), .A2(n6), .ZN(n2) );
  NAND2_X1 U14 ( .A1(port1[30]), .A2(n7), .ZN(n3) );
  INV_X1 U15 ( .A(n33), .ZN(N29) );
  AOI22_X1 U16 ( .A1(port0[27]), .A2(n6), .B1(port1[27]), .B2(n11), .ZN(n33)
         );
  AOI22_X1 U17 ( .A1(port0[26]), .A2(n6), .B1(port1[26]), .B2(n8), .ZN(n32) );
  INV_X1 U18 ( .A(n31), .ZN(N27) );
  AOI22_X1 U19 ( .A1(port0[25]), .A2(n6), .B1(port1[25]), .B2(n9), .ZN(n31) );
  INV_X1 U20 ( .A(n44), .ZN(N31) );
  AOI22_X1 U21 ( .A1(port0[29]), .A2(n6), .B1(port1[29]), .B2(n10), .ZN(n44)
         );
  AOI22_X1 U22 ( .A1(port0[28]), .A2(n6), .B1(port1[28]), .B2(n7), .ZN(n42) );
  AOI22_X1 U23 ( .A1(port0[18]), .A2(n6), .B1(port1[18]), .B2(n11), .ZN(n24)
         );
  INV_X1 U24 ( .A(n30), .ZN(N26) );
  AOI22_X1 U25 ( .A1(port0[24]), .A2(n6), .B1(port1[24]), .B2(n8), .ZN(n30) );
  INV_X1 U26 ( .A(n20), .ZN(N17) );
  AOI22_X1 U27 ( .A1(port0[15]), .A2(n6), .B1(port1[15]), .B2(n9), .ZN(n20) );
  INV_X1 U28 ( .A(n21), .ZN(N18) );
  AOI22_X1 U29 ( .A1(port0[16]), .A2(n6), .B1(port1[16]), .B2(n9), .ZN(n21) );
  AOI22_X1 U30 ( .A1(port0[20]), .A2(n6), .B1(port1[20]), .B2(n10), .ZN(n26)
         );
  AOI22_X1 U32 ( .A1(port0[17]), .A2(n6), .B1(port1[17]), .B2(n9), .ZN(n22) );
  INV_X1 U33 ( .A(n19), .ZN(N16) );
  AOI22_X1 U34 ( .A1(port0[14]), .A2(n6), .B1(port1[14]), .B2(n10), .ZN(n19)
         );
  AOI22_X1 U35 ( .A1(port0[19]), .A2(n6), .B1(port1[19]), .B2(n9), .ZN(n25) );
  INV_X1 U36 ( .A(n18), .ZN(N15) );
  AOI22_X1 U37 ( .A1(port0[13]), .A2(n6), .B1(port1[13]), .B2(n10), .ZN(n18)
         );
  INV_X1 U38 ( .A(n15), .ZN(N12) );
  AOI22_X1 U39 ( .A1(port0[10]), .A2(n6), .B1(port1[10]), .B2(n11), .ZN(n15)
         );
  AOI22_X1 U40 ( .A1(port0[22]), .A2(n6), .B1(port1[22]), .B2(n8), .ZN(n28) );
  AOI22_X1 U41 ( .A1(port0[23]), .A2(n6), .B1(port1[23]), .B2(n8), .ZN(n29) );
  AOI22_X1 U42 ( .A1(port0[21]), .A2(n6), .B1(port1[21]), .B2(n8), .ZN(n27) );
  INV_X1 U43 ( .A(n17), .ZN(N14) );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n6), .B1(port1[12]), .B2(n10), .ZN(n17)
         );
  INV_X1 U45 ( .A(n16), .ZN(N13) );
  AOI22_X1 U46 ( .A1(port0[11]), .A2(n6), .B1(port1[11]), .B2(n10), .ZN(n16)
         );
  INV_X1 U47 ( .A(n14), .ZN(N11) );
  AOI22_X1 U48 ( .A1(port0[9]), .A2(n6), .B1(port1[9]), .B2(n11), .ZN(n14) );
  INV_X1 U49 ( .A(n47), .ZN(N5) );
  AOI22_X1 U50 ( .A1(port0[3]), .A2(n6), .B1(port1[3]), .B2(n11), .ZN(n47) );
  INV_X1 U51 ( .A(n50), .ZN(N8) );
  AOI22_X1 U52 ( .A1(port0[6]), .A2(n6), .B1(port1[6]), .B2(n11), .ZN(n50) );
  INV_X1 U53 ( .A(n35), .ZN(N3) );
  AOI22_X1 U54 ( .A1(port0[1]), .A2(n6), .B1(port1[1]), .B2(n9), .ZN(n35) );
  INV_X1 U55 ( .A(n23), .ZN(N2) );
  AOI22_X1 U56 ( .A1(port0[0]), .A2(n6), .B1(port1[0]), .B2(n9), .ZN(n23) );
  INV_X1 U57 ( .A(n13), .ZN(N10) );
  AOI22_X1 U58 ( .A1(port0[8]), .A2(n6), .B1(port1[8]), .B2(n11), .ZN(n13) );
  INV_X1 U59 ( .A(n49), .ZN(N7) );
  AOI22_X1 U60 ( .A1(port0[5]), .A2(n6), .B1(port1[5]), .B2(n11), .ZN(n49) );
  INV_X1 U61 ( .A(n48), .ZN(N6) );
  AOI22_X1 U62 ( .A1(port0[4]), .A2(n6), .B1(port1[4]), .B2(n11), .ZN(n48) );
  INV_X1 U63 ( .A(n46), .ZN(N4) );
  AOI22_X1 U64 ( .A1(port0[2]), .A2(n6), .B1(port1[2]), .B2(n7), .ZN(n46) );
  INV_X1 U65 ( .A(n51), .ZN(N9) );
  AOI22_X1 U66 ( .A1(port0[7]), .A2(n6), .B1(n11), .B2(port1[7]), .ZN(n51) );
  CLKBUF_X1 U67 ( .A(n10), .Z(n8) );
  CLKBUF_X1 U68 ( .A(n11), .Z(n9) );
  CLKBUF_X1 U69 ( .A(n5), .Z(n10) );
  CLKBUF_X1 U70 ( .A(n5), .Z(n11) );
  BUF_X1 U71 ( .A(sel), .Z(n5) );
  CLKBUF_X1 U72 ( .A(sel), .Z(n4) );
  INV_X1 U73 ( .A(n45), .ZN(N33) );
  AOI22_X1 U74 ( .A1(port0[31]), .A2(n6), .B1(port1[31]), .B2(n7), .ZN(n45) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_78 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n5), .Z(n14) );
  BUF_X1 U5 ( .A(n4), .Z(n11) );
  BUF_X1 U6 ( .A(n4), .Z(n10) );
  BUF_X1 U7 ( .A(n6), .Z(n17) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n61), .ZN(N6) );
  INV_X1 U16 ( .A(n60), .ZN(N5) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  INV_X1 U18 ( .A(n28), .ZN(N2) );
  INV_X1 U19 ( .A(n54), .ZN(N3) );
  INV_X1 U20 ( .A(n62), .ZN(N7) );
  INV_X1 U21 ( .A(n64), .ZN(N9) );
  INV_X1 U22 ( .A(n63), .ZN(N8) );
  INV_X1 U23 ( .A(n58), .ZN(N33) );
  INV_X1 U24 ( .A(n57), .ZN(N32) );
  INV_X1 U25 ( .A(n26), .ZN(N18) );
  INV_X1 U26 ( .A(n31), .ZN(N22) );
  INV_X1 U27 ( .A(n32), .ZN(N23) );
  INV_X1 U28 ( .A(n33), .ZN(N24) );
  INV_X1 U29 ( .A(n35), .ZN(N25) );
  INV_X1 U30 ( .A(n50), .ZN(N26) );
  INV_X1 U31 ( .A(n51), .ZN(N27) );
  INV_X1 U32 ( .A(n52), .ZN(N28) );
  INV_X1 U33 ( .A(n53), .ZN(N29) );
  INV_X1 U34 ( .A(n55), .ZN(N30) );
  INV_X1 U35 ( .A(n56), .ZN(N31) );
  INV_X1 U36 ( .A(n27), .ZN(N19) );
  INV_X1 U37 ( .A(n23), .ZN(N15) );
  INV_X1 U38 ( .A(n22), .ZN(N14) );
  INV_X1 U39 ( .A(n24), .ZN(N16) );
  INV_X1 U40 ( .A(n25), .ZN(N17) );
  INV_X1 U41 ( .A(n21), .ZN(N13) );
  INV_X1 U42 ( .A(n29), .ZN(N20) );
  INV_X1 U43 ( .A(n30), .ZN(N21) );
  INV_X1 U44 ( .A(n20), .ZN(N12) );
  INV_X1 U45 ( .A(n19), .ZN(N11) );
  INV_X1 U46 ( .A(n18), .ZN(N10) );
  AOI22_X1 U47 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U48 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U49 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U50 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U51 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U52 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U53 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U54 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U55 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U56 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U57 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U58 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U59 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U60 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U61 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U62 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U63 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U64 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U65 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U66 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_77 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n5), .Z(n14) );
  BUF_X1 U5 ( .A(n4), .Z(n11) );
  BUF_X1 U6 ( .A(n4), .Z(n10) );
  BUF_X1 U7 ( .A(n6), .Z(n17) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n61), .ZN(N6) );
  INV_X1 U16 ( .A(n60), .ZN(N5) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  INV_X1 U18 ( .A(n28), .ZN(N2) );
  INV_X1 U19 ( .A(n54), .ZN(N3) );
  INV_X1 U20 ( .A(n62), .ZN(N7) );
  INV_X1 U21 ( .A(n64), .ZN(N9) );
  INV_X1 U22 ( .A(n63), .ZN(N8) );
  INV_X1 U23 ( .A(n58), .ZN(N33) );
  INV_X1 U24 ( .A(n57), .ZN(N32) );
  INV_X1 U25 ( .A(n30), .ZN(N21) );
  INV_X1 U26 ( .A(n25), .ZN(N17) );
  INV_X1 U27 ( .A(n26), .ZN(N18) );
  INV_X1 U28 ( .A(n31), .ZN(N22) );
  INV_X1 U29 ( .A(n32), .ZN(N23) );
  INV_X1 U30 ( .A(n33), .ZN(N24) );
  INV_X1 U31 ( .A(n35), .ZN(N25) );
  INV_X1 U32 ( .A(n50), .ZN(N26) );
  INV_X1 U33 ( .A(n51), .ZN(N27) );
  INV_X1 U34 ( .A(n52), .ZN(N28) );
  INV_X1 U35 ( .A(n53), .ZN(N29) );
  INV_X1 U36 ( .A(n55), .ZN(N30) );
  INV_X1 U37 ( .A(n56), .ZN(N31) );
  INV_X1 U38 ( .A(n27), .ZN(N19) );
  INV_X1 U39 ( .A(n23), .ZN(N15) );
  INV_X1 U40 ( .A(n22), .ZN(N14) );
  INV_X1 U41 ( .A(n24), .ZN(N16) );
  INV_X1 U42 ( .A(n21), .ZN(N13) );
  INV_X1 U43 ( .A(n29), .ZN(N20) );
  INV_X1 U44 ( .A(n20), .ZN(N12) );
  INV_X1 U45 ( .A(n19), .ZN(N11) );
  INV_X1 U46 ( .A(n18), .ZN(N10) );
  AOI22_X1 U47 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U48 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U49 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U50 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U51 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U52 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U53 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U54 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U55 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U56 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U57 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U58 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U59 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U60 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U61 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U62 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U63 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U64 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U65 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U66 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_75 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n5), .Z(n14) );
  BUF_X1 U5 ( .A(n4), .Z(n11) );
  BUF_X1 U6 ( .A(n4), .Z(n10) );
  BUF_X1 U7 ( .A(n6), .Z(n17) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n59), .ZN(N4) );
  AOI22_X1 U16 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U17 ( .A(n61), .ZN(N6) );
  AOI22_X1 U18 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U19 ( .A(n60), .ZN(N5) );
  AOI22_X1 U20 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U21 ( .A(n28), .ZN(N2) );
  AOI22_X1 U22 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U23 ( .A(n54), .ZN(N3) );
  AOI22_X1 U24 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U25 ( .A(n27), .ZN(N19) );
  AOI22_X1 U26 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U27 ( .A(n20), .ZN(N12) );
  AOI22_X1 U28 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U29 ( .A(n29), .ZN(N20) );
  AOI22_X1 U30 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U31 ( .A(n31), .ZN(N22) );
  AOI22_X1 U32 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U33 ( .A(n32), .ZN(N23) );
  AOI22_X1 U34 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U35 ( .A(n33), .ZN(N24) );
  AOI22_X1 U36 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U37 ( .A(n35), .ZN(N25) );
  AOI22_X1 U38 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U39 ( .A(n50), .ZN(N26) );
  AOI22_X1 U40 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U41 ( .A(n51), .ZN(N27) );
  AOI22_X1 U42 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U43 ( .A(n52), .ZN(N28) );
  AOI22_X1 U44 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U45 ( .A(n53), .ZN(N29) );
  AOI22_X1 U46 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U47 ( .A(n55), .ZN(N30) );
  AOI22_X1 U48 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U49 ( .A(n56), .ZN(N31) );
  AOI22_X1 U50 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U51 ( .A(n62), .ZN(N7) );
  AOI22_X1 U52 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U53 ( .A(n64), .ZN(N9) );
  AOI22_X1 U54 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U55 ( .A(n63), .ZN(N8) );
  AOI22_X1 U56 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U57 ( .A(n58), .ZN(N33) );
  AOI22_X1 U58 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U59 ( .A(n57), .ZN(N32) );
  AOI22_X1 U60 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U61 ( .A(n23), .ZN(N15) );
  AOI22_X1 U62 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U63 ( .A(n22), .ZN(N14) );
  AOI22_X1 U64 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U65 ( .A(n24), .ZN(N16) );
  AOI22_X1 U66 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U67 ( .A(n19), .ZN(N11) );
  AOI22_X1 U68 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U69 ( .A(n25), .ZN(N17) );
  AOI22_X1 U70 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U71 ( .A(n18), .ZN(N10) );
  AOI22_X1 U72 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U73 ( .A(n21), .ZN(N13) );
  AOI22_X1 U74 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U75 ( .A(n26), .ZN(N18) );
  AOI22_X1 U76 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U77 ( .A(n30), .ZN(N21) );
  AOI22_X1 U78 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_74 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n5), .Z(n14) );
  BUF_X1 U5 ( .A(n4), .Z(n11) );
  BUF_X1 U6 ( .A(n4), .Z(n10) );
  BUF_X1 U7 ( .A(n6), .Z(n17) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n28), .ZN(N2) );
  AOI22_X1 U16 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U17 ( .A(n54), .ZN(N3) );
  AOI22_X1 U18 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U19 ( .A(n61), .ZN(N6) );
  AOI22_X1 U20 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U21 ( .A(n60), .ZN(N5) );
  AOI22_X1 U22 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U23 ( .A(n59), .ZN(N4) );
  AOI22_X1 U24 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U25 ( .A(n62), .ZN(N7) );
  AOI22_X1 U26 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U27 ( .A(n64), .ZN(N9) );
  AOI22_X1 U28 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U29 ( .A(n57), .ZN(N32) );
  AOI22_X1 U30 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U31 ( .A(n25), .ZN(N17) );
  AOI22_X1 U32 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U33 ( .A(n26), .ZN(N18) );
  AOI22_X1 U34 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U35 ( .A(n33), .ZN(N24) );
  AOI22_X1 U36 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U37 ( .A(n35), .ZN(N25) );
  AOI22_X1 U38 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U39 ( .A(n50), .ZN(N26) );
  AOI22_X1 U40 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U41 ( .A(n51), .ZN(N27) );
  AOI22_X1 U42 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U43 ( .A(n52), .ZN(N28) );
  AOI22_X1 U44 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U45 ( .A(n53), .ZN(N29) );
  AOI22_X1 U46 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U47 ( .A(n55), .ZN(N30) );
  AOI22_X1 U48 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U49 ( .A(n56), .ZN(N31) );
  AOI22_X1 U50 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U51 ( .A(n63), .ZN(N8) );
  AOI22_X1 U52 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U53 ( .A(n58), .ZN(N33) );
  AOI22_X1 U54 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U55 ( .A(n27), .ZN(N19) );
  AOI22_X1 U56 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U57 ( .A(n20), .ZN(N12) );
  AOI22_X1 U58 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U59 ( .A(n23), .ZN(N15) );
  AOI22_X1 U60 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U61 ( .A(n22), .ZN(N14) );
  AOI22_X1 U62 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U63 ( .A(n24), .ZN(N16) );
  AOI22_X1 U64 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U65 ( .A(n19), .ZN(N11) );
  AOI22_X1 U66 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U67 ( .A(n18), .ZN(N10) );
  AOI22_X1 U68 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U69 ( .A(n21), .ZN(N13) );
  AOI22_X1 U70 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U71 ( .A(n29), .ZN(N20) );
  AOI22_X1 U72 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U73 ( .A(n30), .ZN(N21) );
  AOI22_X1 U74 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U75 ( .A(n31), .ZN(N22) );
  AOI22_X1 U76 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U77 ( .A(n32), .ZN(N23) );
  AOI22_X1 U78 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_73 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n8) );
  INV_X1 U2 ( .A(n17), .ZN(n7) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n4), .Z(n11) );
  BUF_X1 U5 ( .A(n4), .Z(n10) );
  BUF_X1 U6 ( .A(n5), .Z(n14) );
  BUF_X1 U7 ( .A(n6), .Z(n17) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n12) );
  BUF_X1 U11 ( .A(n5), .Z(n13) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n4) );
  BUF_X1 U14 ( .A(sel), .Z(n5) );
  INV_X1 U15 ( .A(n61), .ZN(N6) );
  AOI22_X1 U16 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U17 ( .A(n60), .ZN(N5) );
  AOI22_X1 U18 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U19 ( .A(n59), .ZN(N4) );
  AOI22_X1 U20 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U21 ( .A(n28), .ZN(N2) );
  AOI22_X1 U22 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U23 ( .A(n54), .ZN(N3) );
  AOI22_X1 U24 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U25 ( .A(n62), .ZN(N7) );
  AOI22_X1 U26 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U27 ( .A(n64), .ZN(N9) );
  AOI22_X1 U28 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U29 ( .A(n63), .ZN(N8) );
  AOI22_X1 U30 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U31 ( .A(n58), .ZN(N33) );
  AOI22_X1 U32 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U33 ( .A(n57), .ZN(N32) );
  AOI22_X1 U34 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U35 ( .A(n29), .ZN(N20) );
  AOI22_X1 U36 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U37 ( .A(n27), .ZN(N19) );
  AOI22_X1 U38 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U39 ( .A(n20), .ZN(N12) );
  AOI22_X1 U40 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U41 ( .A(n23), .ZN(N15) );
  AOI22_X1 U42 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U43 ( .A(n22), .ZN(N14) );
  AOI22_X1 U44 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U45 ( .A(n24), .ZN(N16) );
  AOI22_X1 U46 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U47 ( .A(n19), .ZN(N11) );
  AOI22_X1 U48 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U49 ( .A(n18), .ZN(N10) );
  AOI22_X1 U50 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U51 ( .A(n21), .ZN(N13) );
  AOI22_X1 U52 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U53 ( .A(n30), .ZN(N21) );
  AOI22_X1 U54 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U55 ( .A(n31), .ZN(N22) );
  AOI22_X1 U56 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U57 ( .A(n32), .ZN(N23) );
  AOI22_X1 U58 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U59 ( .A(n25), .ZN(N17) );
  AOI22_X1 U60 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U61 ( .A(n26), .ZN(N18) );
  AOI22_X1 U62 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U63 ( .A(n33), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U65 ( .A(n35), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U67 ( .A(n50), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U69 ( .A(n51), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U71 ( .A(n52), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U73 ( .A(n53), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U75 ( .A(n55), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_71 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n5), .Z(n14) );
  BUF_X1 U5 ( .A(n4), .Z(n11) );
  BUF_X1 U6 ( .A(n4), .Z(n10) );
  BUF_X1 U7 ( .A(n6), .Z(n17) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n61), .ZN(N6) );
  INV_X1 U16 ( .A(n60), .ZN(N5) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  INV_X1 U18 ( .A(n54), .ZN(N3) );
  INV_X1 U19 ( .A(n62), .ZN(N7) );
  INV_X1 U20 ( .A(n64), .ZN(N9) );
  INV_X1 U21 ( .A(n63), .ZN(N8) );
  INV_X1 U22 ( .A(n58), .ZN(N33) );
  INV_X1 U23 ( .A(n57), .ZN(N32) );
  INV_X1 U24 ( .A(n22), .ZN(N14) );
  INV_X1 U25 ( .A(n26), .ZN(N18) );
  INV_X1 U26 ( .A(n31), .ZN(N22) );
  INV_X1 U27 ( .A(n32), .ZN(N23) );
  INV_X1 U28 ( .A(n33), .ZN(N24) );
  INV_X1 U29 ( .A(n35), .ZN(N25) );
  INV_X1 U30 ( .A(n50), .ZN(N26) );
  INV_X1 U31 ( .A(n51), .ZN(N27) );
  INV_X1 U32 ( .A(n52), .ZN(N28) );
  INV_X1 U33 ( .A(n53), .ZN(N29) );
  INV_X1 U34 ( .A(n55), .ZN(N30) );
  INV_X1 U35 ( .A(n56), .ZN(N31) );
  INV_X1 U36 ( .A(n27), .ZN(N19) );
  INV_X1 U37 ( .A(n23), .ZN(N15) );
  INV_X1 U38 ( .A(n24), .ZN(N16) );
  INV_X1 U39 ( .A(n25), .ZN(N17) );
  INV_X1 U40 ( .A(n21), .ZN(N13) );
  INV_X1 U41 ( .A(n29), .ZN(N20) );
  INV_X1 U42 ( .A(n30), .ZN(N21) );
  INV_X1 U43 ( .A(n20), .ZN(N12) );
  INV_X1 U44 ( .A(n19), .ZN(N11) );
  INV_X1 U45 ( .A(n18), .ZN(N10) );
  AOI22_X1 U46 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U47 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U48 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U49 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U50 ( .A(n28), .ZN(N2) );
  AOI22_X1 U51 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U52 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U53 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U54 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U55 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U56 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U57 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U58 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U59 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U60 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U61 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U62 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U63 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U64 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U65 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U66 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_70 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n5), .Z(n14) );
  BUF_X1 U5 ( .A(n4), .Z(n11) );
  BUF_X1 U6 ( .A(n4), .Z(n10) );
  BUF_X1 U7 ( .A(n6), .Z(n17) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n61), .ZN(N6) );
  INV_X1 U16 ( .A(n60), .ZN(N5) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  INV_X1 U18 ( .A(n54), .ZN(N3) );
  INV_X1 U19 ( .A(n62), .ZN(N7) );
  INV_X1 U20 ( .A(n64), .ZN(N9) );
  INV_X1 U21 ( .A(n63), .ZN(N8) );
  INV_X1 U22 ( .A(n58), .ZN(N33) );
  INV_X1 U23 ( .A(n57), .ZN(N32) );
  INV_X1 U24 ( .A(n22), .ZN(N14) );
  INV_X1 U25 ( .A(n26), .ZN(N18) );
  INV_X1 U26 ( .A(n31), .ZN(N22) );
  INV_X1 U27 ( .A(n32), .ZN(N23) );
  INV_X1 U28 ( .A(n33), .ZN(N24) );
  INV_X1 U29 ( .A(n35), .ZN(N25) );
  INV_X1 U30 ( .A(n50), .ZN(N26) );
  INV_X1 U31 ( .A(n51), .ZN(N27) );
  INV_X1 U32 ( .A(n52), .ZN(N28) );
  INV_X1 U33 ( .A(n53), .ZN(N29) );
  INV_X1 U34 ( .A(n55), .ZN(N30) );
  INV_X1 U35 ( .A(n56), .ZN(N31) );
  INV_X1 U36 ( .A(n27), .ZN(N19) );
  INV_X1 U37 ( .A(n23), .ZN(N15) );
  INV_X1 U38 ( .A(n24), .ZN(N16) );
  INV_X1 U39 ( .A(n25), .ZN(N17) );
  INV_X1 U40 ( .A(n21), .ZN(N13) );
  INV_X1 U41 ( .A(n29), .ZN(N20) );
  INV_X1 U42 ( .A(n30), .ZN(N21) );
  INV_X1 U43 ( .A(n20), .ZN(N12) );
  INV_X1 U44 ( .A(n19), .ZN(N11) );
  INV_X1 U45 ( .A(n18), .ZN(N10) );
  AOI22_X1 U46 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U47 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U48 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U49 ( .A(n28), .ZN(N2) );
  AOI22_X1 U50 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U51 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U52 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U53 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U54 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U55 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U56 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U57 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U58 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U59 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U60 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U61 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U62 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U63 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U64 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U65 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U66 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_69 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n8) );
  INV_X1 U2 ( .A(n17), .ZN(n7) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n4), .Z(n11) );
  BUF_X1 U5 ( .A(n4), .Z(n10) );
  BUF_X1 U6 ( .A(n5), .Z(n14) );
  BUF_X1 U7 ( .A(n6), .Z(n17) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n61), .ZN(N6) );
  INV_X1 U16 ( .A(n60), .ZN(N5) );
  INV_X1 U17 ( .A(n59), .ZN(N4) );
  INV_X1 U18 ( .A(n54), .ZN(N3) );
  INV_X1 U19 ( .A(n62), .ZN(N7) );
  INV_X1 U20 ( .A(n58), .ZN(N33) );
  INV_X1 U21 ( .A(n57), .ZN(N32) );
  INV_X1 U22 ( .A(n24), .ZN(N16) );
  INV_X1 U23 ( .A(n21), .ZN(N13) );
  INV_X1 U24 ( .A(n30), .ZN(N21) );
  INV_X1 U25 ( .A(n31), .ZN(N22) );
  INV_X1 U26 ( .A(n32), .ZN(N23) );
  INV_X1 U27 ( .A(n64), .ZN(N9) );
  INV_X1 U28 ( .A(n63), .ZN(N8) );
  INV_X1 U29 ( .A(n25), .ZN(N17) );
  INV_X1 U30 ( .A(n26), .ZN(N18) );
  INV_X1 U31 ( .A(n33), .ZN(N24) );
  INV_X1 U32 ( .A(n35), .ZN(N25) );
  INV_X1 U33 ( .A(n50), .ZN(N26) );
  INV_X1 U34 ( .A(n51), .ZN(N27) );
  INV_X1 U35 ( .A(n52), .ZN(N28) );
  INV_X1 U36 ( .A(n53), .ZN(N29) );
  INV_X1 U37 ( .A(n55), .ZN(N30) );
  INV_X1 U38 ( .A(n56), .ZN(N31) );
  INV_X1 U39 ( .A(n29), .ZN(N20) );
  INV_X1 U40 ( .A(n27), .ZN(N19) );
  INV_X1 U41 ( .A(n23), .ZN(N15) );
  INV_X1 U42 ( .A(n22), .ZN(N14) );
  INV_X1 U43 ( .A(n20), .ZN(N12) );
  INV_X1 U44 ( .A(n19), .ZN(N11) );
  INV_X1 U45 ( .A(n18), .ZN(N10) );
  AOI22_X1 U46 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U47 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U48 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U49 ( .A(n28), .ZN(N2) );
  AOI22_X1 U50 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U51 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U52 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U53 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U54 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U55 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U56 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U57 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U58 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U59 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U60 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U61 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U62 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U63 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U64 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U65 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U66 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_67 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n5), .Z(n14) );
  BUF_X1 U5 ( .A(n4), .Z(n11) );
  BUF_X1 U6 ( .A(n4), .Z(n10) );
  BUF_X1 U7 ( .A(n6), .Z(n17) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n28), .ZN(N2) );
  INV_X1 U16 ( .A(n59), .ZN(N4) );
  AOI22_X1 U17 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U18 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U19 ( .A(n61), .ZN(N6) );
  AOI22_X1 U20 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U21 ( .A(n60), .ZN(N5) );
  AOI22_X1 U22 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U23 ( .A(n54), .ZN(N3) );
  AOI22_X1 U24 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U25 ( .A(n27), .ZN(N19) );
  AOI22_X1 U26 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U27 ( .A(n20), .ZN(N12) );
  AOI22_X1 U28 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U29 ( .A(n29), .ZN(N20) );
  AOI22_X1 U30 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U31 ( .A(n31), .ZN(N22) );
  AOI22_X1 U32 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U33 ( .A(n32), .ZN(N23) );
  AOI22_X1 U34 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U35 ( .A(n33), .ZN(N24) );
  AOI22_X1 U36 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U37 ( .A(n35), .ZN(N25) );
  AOI22_X1 U38 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U39 ( .A(n50), .ZN(N26) );
  AOI22_X1 U40 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U41 ( .A(n51), .ZN(N27) );
  AOI22_X1 U42 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U43 ( .A(n52), .ZN(N28) );
  AOI22_X1 U44 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U45 ( .A(n53), .ZN(N29) );
  AOI22_X1 U46 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U47 ( .A(n55), .ZN(N30) );
  AOI22_X1 U48 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U49 ( .A(n56), .ZN(N31) );
  AOI22_X1 U50 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U51 ( .A(n62), .ZN(N7) );
  AOI22_X1 U52 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U53 ( .A(n64), .ZN(N9) );
  AOI22_X1 U54 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U55 ( .A(n63), .ZN(N8) );
  AOI22_X1 U56 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U57 ( .A(n58), .ZN(N33) );
  AOI22_X1 U58 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U59 ( .A(n57), .ZN(N32) );
  AOI22_X1 U60 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U61 ( .A(n23), .ZN(N15) );
  AOI22_X1 U62 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U63 ( .A(n22), .ZN(N14) );
  AOI22_X1 U64 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U65 ( .A(n24), .ZN(N16) );
  AOI22_X1 U66 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U67 ( .A(n19), .ZN(N11) );
  AOI22_X1 U68 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U69 ( .A(n25), .ZN(N17) );
  AOI22_X1 U70 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U71 ( .A(n18), .ZN(N10) );
  AOI22_X1 U72 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U73 ( .A(n21), .ZN(N13) );
  AOI22_X1 U74 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U75 ( .A(n26), .ZN(N18) );
  AOI22_X1 U76 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U77 ( .A(n30), .ZN(N21) );
  AOI22_X1 U78 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_66 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n5), .Z(n14) );
  BUF_X1 U5 ( .A(n4), .Z(n11) );
  BUF_X1 U6 ( .A(n4), .Z(n10) );
  BUF_X1 U7 ( .A(n6), .Z(n17) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n28), .ZN(N2) );
  AOI22_X1 U16 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U17 ( .A(n54), .ZN(N3) );
  AOI22_X1 U18 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U19 ( .A(n61), .ZN(N6) );
  AOI22_X1 U20 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U21 ( .A(n60), .ZN(N5) );
  AOI22_X1 U22 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U23 ( .A(n59), .ZN(N4) );
  AOI22_X1 U24 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U25 ( .A(n62), .ZN(N7) );
  AOI22_X1 U26 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U27 ( .A(n57), .ZN(N32) );
  AOI22_X1 U28 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U29 ( .A(n22), .ZN(N14) );
  AOI22_X1 U30 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U31 ( .A(n25), .ZN(N17) );
  AOI22_X1 U32 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U33 ( .A(n26), .ZN(N18) );
  AOI22_X1 U34 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U35 ( .A(n50), .ZN(N26) );
  AOI22_X1 U36 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U37 ( .A(n51), .ZN(N27) );
  AOI22_X1 U38 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U39 ( .A(n52), .ZN(N28) );
  AOI22_X1 U40 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U41 ( .A(n53), .ZN(N29) );
  AOI22_X1 U42 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U43 ( .A(n55), .ZN(N30) );
  AOI22_X1 U44 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U45 ( .A(n56), .ZN(N31) );
  AOI22_X1 U46 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U47 ( .A(n64), .ZN(N9) );
  AOI22_X1 U48 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U49 ( .A(n63), .ZN(N8) );
  AOI22_X1 U50 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U51 ( .A(n58), .ZN(N33) );
  AOI22_X1 U52 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U53 ( .A(n29), .ZN(N20) );
  AOI22_X1 U54 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U55 ( .A(n27), .ZN(N19) );
  AOI22_X1 U56 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U57 ( .A(n20), .ZN(N12) );
  AOI22_X1 U58 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U59 ( .A(n23), .ZN(N15) );
  AOI22_X1 U60 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U61 ( .A(n24), .ZN(N16) );
  AOI22_X1 U62 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U63 ( .A(n19), .ZN(N11) );
  AOI22_X1 U64 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U65 ( .A(n18), .ZN(N10) );
  AOI22_X1 U66 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U67 ( .A(n21), .ZN(N13) );
  AOI22_X1 U68 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U69 ( .A(n30), .ZN(N21) );
  AOI22_X1 U70 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U71 ( .A(n31), .ZN(N22) );
  AOI22_X1 U72 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U73 ( .A(n32), .ZN(N23) );
  AOI22_X1 U74 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U75 ( .A(n33), .ZN(N24) );
  AOI22_X1 U76 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U77 ( .A(n35), .ZN(N25) );
  AOI22_X1 U78 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_65 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n5), .Z(n14) );
  BUF_X1 U5 ( .A(n4), .Z(n11) );
  BUF_X1 U6 ( .A(n4), .Z(n10) );
  BUF_X1 U7 ( .A(n6), .Z(n17) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n12) );
  BUF_X1 U11 ( .A(n5), .Z(n13) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n28), .ZN(N2) );
  INV_X1 U16 ( .A(n61), .ZN(N6) );
  AOI22_X1 U17 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U18 ( .A(n60), .ZN(N5) );
  AOI22_X1 U19 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U20 ( .A(n59), .ZN(N4) );
  AOI22_X1 U21 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U22 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U23 ( .A(n54), .ZN(N3) );
  AOI22_X1 U24 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U25 ( .A(n62), .ZN(N7) );
  AOI22_X1 U26 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U27 ( .A(n64), .ZN(N9) );
  AOI22_X1 U28 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U29 ( .A(n63), .ZN(N8) );
  AOI22_X1 U30 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U31 ( .A(n58), .ZN(N33) );
  AOI22_X1 U32 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U33 ( .A(n57), .ZN(N32) );
  AOI22_X1 U34 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U35 ( .A(n29), .ZN(N20) );
  AOI22_X1 U36 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U37 ( .A(n27), .ZN(N19) );
  AOI22_X1 U38 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U39 ( .A(n20), .ZN(N12) );
  AOI22_X1 U40 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U41 ( .A(n23), .ZN(N15) );
  AOI22_X1 U42 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U43 ( .A(n24), .ZN(N16) );
  AOI22_X1 U44 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U45 ( .A(n22), .ZN(N14) );
  AOI22_X1 U46 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U47 ( .A(n19), .ZN(N11) );
  AOI22_X1 U48 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U49 ( .A(n25), .ZN(N17) );
  AOI22_X1 U50 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U51 ( .A(n18), .ZN(N10) );
  AOI22_X1 U52 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U53 ( .A(n21), .ZN(N13) );
  AOI22_X1 U54 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U55 ( .A(n30), .ZN(N21) );
  AOI22_X1 U56 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U57 ( .A(n31), .ZN(N22) );
  AOI22_X1 U58 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U59 ( .A(n32), .ZN(N23) );
  AOI22_X1 U60 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U61 ( .A(n33), .ZN(N24) );
  AOI22_X1 U62 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U63 ( .A(n35), .ZN(N25) );
  AOI22_X1 U64 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U65 ( .A(n26), .ZN(N18) );
  AOI22_X1 U66 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U67 ( .A(n50), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U69 ( .A(n51), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U71 ( .A(n52), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U73 ( .A(n53), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U75 ( .A(n55), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_64 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n5), .Z(n14) );
  BUF_X1 U5 ( .A(n4), .Z(n11) );
  BUF_X1 U6 ( .A(n4), .Z(n10) );
  BUF_X1 U7 ( .A(n6), .Z(n17) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n28), .ZN(N2) );
  INV_X1 U16 ( .A(n61), .ZN(N6) );
  INV_X1 U17 ( .A(n60), .ZN(N5) );
  AOI22_X1 U18 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U19 ( .A(n59), .ZN(N4) );
  AOI22_X1 U20 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U21 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U22 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U23 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U24 ( .A(n54), .ZN(N3) );
  INV_X1 U25 ( .A(n62), .ZN(N7) );
  AOI22_X1 U26 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U27 ( .A(n64), .ZN(N9) );
  AOI22_X1 U28 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U29 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U30 ( .A(n63), .ZN(N8) );
  AOI22_X1 U31 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U32 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U33 ( .A(n58), .ZN(N33) );
  INV_X1 U34 ( .A(n57), .ZN(N32) );
  INV_X1 U35 ( .A(n29), .ZN(N20) );
  AOI22_X1 U36 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U37 ( .A(n27), .ZN(N19) );
  INV_X1 U38 ( .A(n20), .ZN(N12) );
  INV_X1 U39 ( .A(n23), .ZN(N15) );
  INV_X1 U40 ( .A(n24), .ZN(N16) );
  INV_X1 U41 ( .A(n22), .ZN(N14) );
  INV_X1 U42 ( .A(n19), .ZN(N11) );
  INV_X1 U43 ( .A(n25), .ZN(N17) );
  AOI22_X1 U44 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U45 ( .A(n18), .ZN(N10) );
  AOI22_X1 U46 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U47 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U48 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U49 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U50 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U51 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U52 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U53 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U54 ( .A(n21), .ZN(N13) );
  AOI22_X1 U55 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U56 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U57 ( .A(n30), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U59 ( .A(n31), .ZN(N22) );
  AOI22_X1 U60 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U61 ( .A(n32), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U63 ( .A(n33), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U65 ( .A(n35), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U67 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U68 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U69 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U70 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U71 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U72 ( .A(n26), .ZN(N18) );
  INV_X1 U73 ( .A(n50), .ZN(N26) );
  INV_X1 U74 ( .A(n51), .ZN(N27) );
  INV_X1 U75 ( .A(n52), .ZN(N28) );
  INV_X1 U76 ( .A(n53), .ZN(N29) );
  INV_X1 U77 ( .A(n55), .ZN(N30) );
  INV_X1 U78 ( .A(n56), .ZN(N31) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_57 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n5), .Z(n14) );
  BUF_X1 U4 ( .A(n4), .Z(n11) );
  BUF_X1 U5 ( .A(n4), .Z(n10) );
  BUF_X1 U6 ( .A(n6), .Z(n17) );
  BUF_X1 U7 ( .A(n4), .Z(n9) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n12) );
  BUF_X1 U11 ( .A(n5), .Z(n13) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n59), .ZN(N4) );
  AOI22_X1 U16 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U17 ( .A(n54), .ZN(N3) );
  AOI22_X1 U18 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U19 ( .A(n61), .ZN(N6) );
  AOI22_X1 U20 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U21 ( .A(n60), .ZN(N5) );
  AOI22_X1 U22 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U23 ( .A(n28), .ZN(N2) );
  AOI22_X1 U24 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U25 ( .A(n62), .ZN(N7) );
  AOI22_X1 U26 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U27 ( .A(n64), .ZN(N9) );
  AOI22_X1 U28 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U29 ( .A(n29), .ZN(N20) );
  AOI22_X1 U30 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U31 ( .A(n27), .ZN(N19) );
  AOI22_X1 U32 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U33 ( .A(n20), .ZN(N12) );
  AOI22_X1 U34 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U35 ( .A(n23), .ZN(N15) );
  AOI22_X1 U36 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U37 ( .A(n22), .ZN(N14) );
  AOI22_X1 U38 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U39 ( .A(n24), .ZN(N16) );
  AOI22_X1 U40 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U41 ( .A(n19), .ZN(N11) );
  AOI22_X1 U42 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U43 ( .A(n18), .ZN(N10) );
  AOI22_X1 U44 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U45 ( .A(n21), .ZN(N13) );
  AOI22_X1 U46 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U47 ( .A(n26), .ZN(N18) );
  AOI22_X1 U48 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  INV_X1 U49 ( .A(n63), .ZN(N8) );
  AOI22_X1 U50 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U51 ( .A(n58), .ZN(N33) );
  AOI22_X1 U52 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U53 ( .A(n57), .ZN(N32) );
  AOI22_X1 U54 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U55 ( .A(n25), .ZN(N17) );
  AOI22_X1 U56 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U57 ( .A(n30), .ZN(N21) );
  AOI22_X1 U58 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U59 ( .A(n31), .ZN(N22) );
  AOI22_X1 U60 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U61 ( .A(n32), .ZN(N23) );
  AOI22_X1 U62 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U63 ( .A(n33), .ZN(N24) );
  AOI22_X1 U64 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U65 ( .A(n35), .ZN(N25) );
  AOI22_X1 U66 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U67 ( .A(n50), .ZN(N26) );
  AOI22_X1 U68 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U69 ( .A(n51), .ZN(N27) );
  AOI22_X1 U70 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U71 ( .A(n52), .ZN(N28) );
  AOI22_X1 U72 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U73 ( .A(n53), .ZN(N29) );
  AOI22_X1 U74 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U75 ( .A(n55), .ZN(N30) );
  AOI22_X1 U76 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U77 ( .A(n56), .ZN(N31) );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_56 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n5), .Z(n14) );
  BUF_X1 U4 ( .A(n4), .Z(n11) );
  BUF_X1 U5 ( .A(n4), .Z(n10) );
  BUF_X1 U6 ( .A(n6), .Z(n17) );
  BUF_X1 U7 ( .A(n4), .Z(n9) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n59), .ZN(N4) );
  INV_X1 U16 ( .A(n54), .ZN(N3) );
  INV_X1 U17 ( .A(n61), .ZN(N6) );
  INV_X1 U18 ( .A(n60), .ZN(N5) );
  INV_X1 U19 ( .A(n28), .ZN(N2) );
  AOI22_X1 U20 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U21 ( .A(n62), .ZN(N7) );
  INV_X1 U22 ( .A(n64), .ZN(N9) );
  INV_X1 U23 ( .A(n29), .ZN(N20) );
  INV_X1 U24 ( .A(n27), .ZN(N19) );
  INV_X1 U25 ( .A(n20), .ZN(N12) );
  INV_X1 U26 ( .A(n23), .ZN(N15) );
  INV_X1 U27 ( .A(n22), .ZN(N14) );
  INV_X1 U28 ( .A(n24), .ZN(N16) );
  INV_X1 U29 ( .A(n19), .ZN(N11) );
  INV_X1 U30 ( .A(n18), .ZN(N10) );
  INV_X1 U31 ( .A(n21), .ZN(N13) );
  INV_X1 U32 ( .A(n26), .ZN(N18) );
  INV_X1 U33 ( .A(n63), .ZN(N8) );
  INV_X1 U34 ( .A(n58), .ZN(N33) );
  INV_X1 U35 ( .A(n57), .ZN(N32) );
  INV_X1 U36 ( .A(n25), .ZN(N17) );
  INV_X1 U37 ( .A(n30), .ZN(N21) );
  INV_X1 U38 ( .A(n31), .ZN(N22) );
  INV_X1 U39 ( .A(n32), .ZN(N23) );
  INV_X1 U40 ( .A(n33), .ZN(N24) );
  INV_X1 U41 ( .A(n35), .ZN(N25) );
  INV_X1 U42 ( .A(n50), .ZN(N26) );
  INV_X1 U43 ( .A(n51), .ZN(N27) );
  INV_X1 U44 ( .A(n52), .ZN(N28) );
  INV_X1 U45 ( .A(n53), .ZN(N29) );
  INV_X1 U46 ( .A(n55), .ZN(N30) );
  INV_X1 U47 ( .A(n56), .ZN(N31) );
  AOI22_X1 U48 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U49 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U50 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U51 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U52 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U53 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U54 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U55 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U56 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  AOI22_X1 U57 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U58 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U59 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U60 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U61 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U62 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U63 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U64 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U65 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U66 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U67 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U68 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U69 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U70 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U71 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U72 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_55 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n8) );
  INV_X1 U2 ( .A(n17), .ZN(n7) );
  INV_X1 U3 ( .A(n61), .ZN(N6) );
  AOI22_X1 U4 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U5 ( .A(n60), .ZN(N5) );
  AOI22_X1 U6 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U7 ( .A(n28), .ZN(N2) );
  AOI22_X1 U8 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  INV_X1 U9 ( .A(n54), .ZN(N3) );
  AOI22_X1 U10 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U11 ( .A(n59), .ZN(N4) );
  AOI22_X1 U12 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U13 ( .A(n64), .ZN(N9) );
  AOI22_X1 U14 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U15 ( .A(n63), .ZN(N8) );
  AOI22_X1 U16 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U17 ( .A(n27), .ZN(N19) );
  AOI22_X1 U18 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U19 ( .A(n23), .ZN(N15) );
  AOI22_X1 U20 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U21 ( .A(n22), .ZN(N14) );
  AOI22_X1 U22 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U23 ( .A(n19), .ZN(N11) );
  AOI22_X1 U24 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U25 ( .A(n25), .ZN(N17) );
  AOI22_X1 U26 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U27 ( .A(n18), .ZN(N10) );
  AOI22_X1 U28 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U29 ( .A(n21), .ZN(N13) );
  AOI22_X1 U30 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U31 ( .A(n26), .ZN(N18) );
  AOI22_X1 U32 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  BUF_X1 U33 ( .A(n4), .Z(n11) );
  BUF_X1 U34 ( .A(n5), .Z(n14) );
  BUF_X1 U35 ( .A(n6), .Z(n17) );
  INV_X1 U36 ( .A(n62), .ZN(N7) );
  AOI22_X1 U37 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U38 ( .A(n58), .ZN(N33) );
  AOI22_X1 U39 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U40 ( .A(n57), .ZN(N32) );
  AOI22_X1 U41 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U42 ( .A(n29), .ZN(N20) );
  AOI22_X1 U43 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U44 ( .A(n24), .ZN(N16) );
  AOI22_X1 U45 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U46 ( .A(n30), .ZN(N21) );
  AOI22_X1 U47 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U48 ( .A(n31), .ZN(N22) );
  AOI22_X1 U49 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U50 ( .A(n32), .ZN(N23) );
  AOI22_X1 U51 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U52 ( .A(n33), .ZN(N24) );
  AOI22_X1 U53 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U54 ( .A(n35), .ZN(N25) );
  AOI22_X1 U55 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U56 ( .A(n50), .ZN(N26) );
  AOI22_X1 U57 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U58 ( .A(n51), .ZN(N27) );
  AOI22_X1 U59 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U60 ( .A(n52), .ZN(N28) );
  AOI22_X1 U61 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U62 ( .A(n53), .ZN(N29) );
  AOI22_X1 U63 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U64 ( .A(n55), .ZN(N30) );
  AOI22_X1 U65 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U66 ( .A(n56), .ZN(N31) );
  AOI22_X1 U67 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  INV_X1 U68 ( .A(n20), .ZN(N12) );
  AOI22_X1 U69 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  BUF_X1 U70 ( .A(n6), .Z(n15) );
  BUF_X1 U71 ( .A(n4), .Z(n10) );
  BUF_X1 U72 ( .A(n4), .Z(n9) );
  BUF_X1 U73 ( .A(n6), .Z(n16) );
  BUF_X1 U74 ( .A(n5), .Z(n12) );
  BUF_X1 U75 ( .A(n5), .Z(n13) );
  BUF_X1 U76 ( .A(sel), .Z(n6) );
  BUF_X1 U77 ( .A(sel), .Z(n4) );
  BUF_X1 U78 ( .A(sel), .Z(n5) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_54 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  INV_X1 U3 ( .A(n61), .ZN(N6) );
  INV_X1 U4 ( .A(n60), .ZN(N5) );
  INV_X1 U5 ( .A(n28), .ZN(N2) );
  INV_X1 U6 ( .A(n54), .ZN(N3) );
  INV_X1 U7 ( .A(n59), .ZN(N4) );
  INV_X1 U8 ( .A(n64), .ZN(N9) );
  INV_X1 U9 ( .A(n63), .ZN(N8) );
  INV_X1 U10 ( .A(n27), .ZN(N19) );
  INV_X1 U11 ( .A(n23), .ZN(N15) );
  INV_X1 U12 ( .A(n22), .ZN(N14) );
  INV_X1 U13 ( .A(n19), .ZN(N11) );
  INV_X1 U14 ( .A(n25), .ZN(N17) );
  INV_X1 U15 ( .A(n18), .ZN(N10) );
  INV_X1 U16 ( .A(n21), .ZN(N13) );
  INV_X1 U17 ( .A(n26), .ZN(N18) );
  BUF_X1 U18 ( .A(n5), .Z(n14) );
  BUF_X1 U19 ( .A(n4), .Z(n11) );
  BUF_X1 U20 ( .A(n6), .Z(n17) );
  INV_X1 U21 ( .A(n62), .ZN(N7) );
  INV_X1 U22 ( .A(n58), .ZN(N33) );
  INV_X1 U23 ( .A(n57), .ZN(N32) );
  INV_X1 U24 ( .A(n29), .ZN(N20) );
  INV_X1 U25 ( .A(n24), .ZN(N16) );
  INV_X1 U26 ( .A(n30), .ZN(N21) );
  INV_X1 U27 ( .A(n31), .ZN(N22) );
  INV_X1 U28 ( .A(n32), .ZN(N23) );
  INV_X1 U29 ( .A(n33), .ZN(N24) );
  INV_X1 U30 ( .A(n35), .ZN(N25) );
  INV_X1 U31 ( .A(n50), .ZN(N26) );
  INV_X1 U32 ( .A(n51), .ZN(N27) );
  INV_X1 U33 ( .A(n52), .ZN(N28) );
  INV_X1 U34 ( .A(n53), .ZN(N29) );
  INV_X1 U35 ( .A(n55), .ZN(N30) );
  INV_X1 U36 ( .A(n56), .ZN(N31) );
  INV_X1 U37 ( .A(n20), .ZN(N12) );
  BUF_X1 U38 ( .A(n4), .Z(n9) );
  BUF_X1 U39 ( .A(n6), .Z(n15) );
  BUF_X1 U40 ( .A(n4), .Z(n10) );
  BUF_X1 U41 ( .A(n6), .Z(n16) );
  BUF_X1 U42 ( .A(n5), .Z(n13) );
  BUF_X1 U43 ( .A(n5), .Z(n12) );
  AOI22_X1 U44 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  AOI22_X1 U45 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  AOI22_X1 U46 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  AOI22_X1 U47 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  AOI22_X1 U48 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  AOI22_X1 U49 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  AOI22_X1 U50 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  AOI22_X1 U51 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  AOI22_X1 U52 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  AOI22_X1 U53 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  AOI22_X1 U54 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  AOI22_X1 U55 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  AOI22_X1 U56 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  AOI22_X1 U57 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  AOI22_X1 U58 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  AOI22_X1 U59 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  AOI22_X1 U60 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  AOI22_X1 U61 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  AOI22_X1 U62 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  BUF_X1 U63 ( .A(sel), .Z(n6) );
  BUF_X1 U64 ( .A(sel), .Z(n5) );
  BUF_X1 U65 ( .A(sel), .Z(n4) );
  AOI22_X1 U66 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  AOI22_X1 U67 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN32_53 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15,
         n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29,
         n30, n31, n32, n33, n35, n50, n51, n52, n53, n54, n55, n56, n57, n58,
         n59, n60, n61, n62, n63, n64;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  INV_X1 U3 ( .A(n28), .ZN(N2) );
  INV_X1 U4 ( .A(n61), .ZN(N6) );
  AOI22_X1 U5 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n61) );
  INV_X1 U6 ( .A(n60), .ZN(N5) );
  AOI22_X1 U7 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n60) );
  INV_X1 U8 ( .A(n59), .ZN(N4) );
  AOI22_X1 U9 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n59) );
  INV_X1 U10 ( .A(n54), .ZN(N3) );
  AOI22_X1 U11 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n54) );
  INV_X1 U12 ( .A(n64), .ZN(N9) );
  AOI22_X1 U13 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n64) );
  INV_X1 U14 ( .A(n63), .ZN(N8) );
  AOI22_X1 U15 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n63) );
  INV_X1 U16 ( .A(n27), .ZN(N19) );
  AOI22_X1 U17 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n27)
         );
  INV_X1 U18 ( .A(n20), .ZN(N12) );
  AOI22_X1 U19 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n20)
         );
  INV_X1 U20 ( .A(n23), .ZN(N15) );
  AOI22_X1 U21 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n23)
         );
  INV_X1 U22 ( .A(n22), .ZN(N14) );
  AOI22_X1 U23 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n22)
         );
  INV_X1 U24 ( .A(n19), .ZN(N11) );
  AOI22_X1 U25 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n19) );
  INV_X1 U26 ( .A(n25), .ZN(N17) );
  AOI22_X1 U27 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n25)
         );
  INV_X1 U28 ( .A(n18), .ZN(N10) );
  AOI22_X1 U29 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n18) );
  INV_X1 U30 ( .A(n21), .ZN(N13) );
  AOI22_X1 U31 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n21)
         );
  INV_X1 U32 ( .A(n26), .ZN(N18) );
  AOI22_X1 U33 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n26)
         );
  BUF_X1 U34 ( .A(n5), .Z(n14) );
  BUF_X1 U35 ( .A(n4), .Z(n11) );
  BUF_X1 U36 ( .A(n6), .Z(n17) );
  INV_X1 U37 ( .A(n62), .ZN(N7) );
  AOI22_X1 U38 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n62) );
  INV_X1 U39 ( .A(n58), .ZN(N33) );
  AOI22_X1 U40 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n58)
         );
  INV_X1 U41 ( .A(n57), .ZN(N32) );
  AOI22_X1 U42 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n57)
         );
  INV_X1 U43 ( .A(n29), .ZN(N20) );
  AOI22_X1 U44 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n29)
         );
  INV_X1 U45 ( .A(n24), .ZN(N16) );
  AOI22_X1 U46 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n24)
         );
  INV_X1 U47 ( .A(n30), .ZN(N21) );
  AOI22_X1 U48 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n30)
         );
  INV_X1 U49 ( .A(n31), .ZN(N22) );
  AOI22_X1 U50 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n31)
         );
  INV_X1 U51 ( .A(n32), .ZN(N23) );
  AOI22_X1 U52 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n32)
         );
  INV_X1 U53 ( .A(n33), .ZN(N24) );
  AOI22_X1 U54 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n33)
         );
  INV_X1 U55 ( .A(n35), .ZN(N25) );
  AOI22_X1 U56 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n35)
         );
  INV_X1 U57 ( .A(n50), .ZN(N26) );
  AOI22_X1 U58 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n50)
         );
  INV_X1 U59 ( .A(n51), .ZN(N27) );
  AOI22_X1 U60 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n51)
         );
  INV_X1 U61 ( .A(n52), .ZN(N28) );
  AOI22_X1 U62 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n52)
         );
  INV_X1 U63 ( .A(n53), .ZN(N29) );
  AOI22_X1 U64 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n53)
         );
  INV_X1 U65 ( .A(n55), .ZN(N30) );
  AOI22_X1 U66 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n55)
         );
  INV_X1 U67 ( .A(n56), .ZN(N31) );
  AOI22_X1 U68 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n56)
         );
  BUF_X1 U69 ( .A(n6), .Z(n15) );
  BUF_X1 U70 ( .A(n4), .Z(n10) );
  BUF_X1 U71 ( .A(n4), .Z(n9) );
  BUF_X1 U72 ( .A(n6), .Z(n16) );
  BUF_X1 U73 ( .A(n5), .Z(n12) );
  BUF_X1 U74 ( .A(n5), .Z(n13) );
  AOI22_X1 U75 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n28) );
  BUF_X1 U76 ( .A(sel), .Z(n6) );
  BUF_X1 U77 ( .A(sel), .Z(n5) );
  BUF_X1 U78 ( .A(sel), .Z(n4) );
endmodule


module NRegister_N32_115 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, net108226, net108227, net108228, net108229,
         net108230, net108231, net108232, net108233, net108234, net108235,
         net108236, net108237, net108238, net108239, net108240, net108241,
         net108242, net108243, net108244, net108245, net108246, net108247,
         net108248, net108249, net108250, net108251, net108252, net108253,
         net108254, net108255, net108256, net108257, n36, n37, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n48), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n50), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n50), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n50), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n49), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n49), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n49), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n48), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n49), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n50), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n48), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n50), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n49), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n48), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n50), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n50), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n50), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n48), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n48), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n48), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n48), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n48), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n48), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n48), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n48), .Q(data_out[0]), 
        .QN(net108226) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n49), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n49), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n49), .Q(n36), .QN(
        net108246) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n49), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n49), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n49), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n49), .QN(net108245) );
  INV_X2 U3 ( .A(net108245), .ZN(data_out[19]) );
  INV_X1 U4 ( .A(n36), .ZN(n37) );
  INV_X2 U5 ( .A(net108246), .ZN(data_out[20]) );
  INV_X1 U6 ( .A(n47), .ZN(n40) );
  INV_X1 U7 ( .A(n47), .ZN(n39) );
  BUF_X1 U8 ( .A(n98), .Z(n43) );
  BUF_X1 U9 ( .A(n98), .Z(n44) );
  BUF_X1 U10 ( .A(n98), .Z(n46) );
  BUF_X1 U11 ( .A(n98), .Z(n41) );
  BUF_X1 U12 ( .A(n98), .Z(n42) );
  BUF_X1 U13 ( .A(n98), .Z(n45) );
  BUF_X1 U14 ( .A(n98), .Z(n47) );
  BUF_X1 U15 ( .A(n3), .Z(n49) );
  BUF_X1 U16 ( .A(n3), .Z(n48) );
  BUF_X1 U17 ( .A(n3), .Z(n50) );
  OAI22_X1 U18 ( .A1(n42), .A2(n91), .B1(net108226), .B2(n40), .ZN(n34) );
  INV_X1 U19 ( .A(data_in[0]), .ZN(n91) );
  OAI22_X1 U20 ( .A1(n42), .A2(n90), .B1(net108227), .B2(n39), .ZN(n33) );
  INV_X1 U21 ( .A(data_in[1]), .ZN(n90) );
  OAI22_X1 U22 ( .A1(n41), .A2(n97), .B1(net108251), .B2(n40), .ZN(n9) );
  INV_X1 U23 ( .A(data_in[25]), .ZN(n97) );
  OAI22_X1 U24 ( .A1(n41), .A2(n96), .B1(net108252), .B2(n39), .ZN(n8) );
  INV_X1 U25 ( .A(data_in[26]), .ZN(n96) );
  OAI22_X1 U26 ( .A1(n41), .A2(n95), .B1(net108253), .B2(n40), .ZN(n7) );
  INV_X1 U27 ( .A(data_in[27]), .ZN(n95) );
  OAI22_X1 U28 ( .A1(n41), .A2(n94), .B1(net108254), .B2(n39), .ZN(n6) );
  INV_X1 U29 ( .A(data_in[28]), .ZN(n94) );
  OAI22_X1 U30 ( .A1(n41), .A2(n93), .B1(net108255), .B2(n40), .ZN(n5) );
  INV_X1 U31 ( .A(data_in[29]), .ZN(n93) );
  OAI22_X1 U32 ( .A1(n42), .A2(n92), .B1(net108256), .B2(n39), .ZN(n4) );
  INV_X1 U33 ( .A(data_in[30]), .ZN(n92) );
  OAI22_X1 U34 ( .A1(n42), .A2(n89), .B1(net108228), .B2(n40), .ZN(n32) );
  INV_X1 U35 ( .A(data_in[2]), .ZN(n89) );
  OAI22_X1 U36 ( .A1(n42), .A2(n88), .B1(net108229), .B2(n40), .ZN(n31) );
  INV_X1 U37 ( .A(data_in[3]), .ZN(n88) );
  OAI22_X1 U38 ( .A1(n43), .A2(n87), .B1(net108230), .B2(n40), .ZN(n30) );
  INV_X1 U39 ( .A(data_in[4]), .ZN(n87) );
  OAI22_X1 U40 ( .A1(n43), .A2(n86), .B1(net108231), .B2(n40), .ZN(n29) );
  INV_X1 U41 ( .A(data_in[5]), .ZN(n86) );
  OAI22_X1 U42 ( .A1(n43), .A2(n85), .B1(net108232), .B2(n40), .ZN(n28) );
  INV_X1 U43 ( .A(data_in[6]), .ZN(n85) );
  OAI22_X1 U44 ( .A1(n43), .A2(n84), .B1(net108233), .B2(n40), .ZN(n27) );
  INV_X1 U45 ( .A(data_in[7]), .ZN(n84) );
  OAI22_X1 U46 ( .A1(n43), .A2(n70), .B1(net108234), .B2(n40), .ZN(n26) );
  INV_X1 U47 ( .A(data_in[8]), .ZN(n70) );
  OAI22_X1 U48 ( .A1(n44), .A2(n67), .B1(net108235), .B2(n40), .ZN(n25) );
  INV_X1 U49 ( .A(data_in[9]), .ZN(n67) );
  OAI22_X1 U50 ( .A1(n44), .A2(n66), .B1(net108236), .B2(n40), .ZN(n24) );
  INV_X1 U51 ( .A(data_in[10]), .ZN(n66) );
  OAI22_X1 U52 ( .A1(n44), .A2(n65), .B1(net108237), .B2(n40), .ZN(n23) );
  INV_X1 U53 ( .A(data_in[11]), .ZN(n65) );
  OAI22_X1 U54 ( .A1(n44), .A2(n64), .B1(net108238), .B2(n40), .ZN(n22) );
  INV_X1 U55 ( .A(data_in[12]), .ZN(n64) );
  OAI22_X1 U56 ( .A1(n44), .A2(n63), .B1(net108239), .B2(n40), .ZN(n21) );
  INV_X1 U57 ( .A(data_in[13]), .ZN(n63) );
  OAI22_X1 U58 ( .A1(n45), .A2(n62), .B1(net108240), .B2(n39), .ZN(n20) );
  INV_X1 U59 ( .A(data_in[14]), .ZN(n62) );
  OAI22_X1 U60 ( .A1(n45), .A2(n60), .B1(net108241), .B2(n39), .ZN(n19) );
  INV_X1 U61 ( .A(data_in[15]), .ZN(n60) );
  OAI22_X1 U62 ( .A1(n45), .A2(n59), .B1(net108242), .B2(n39), .ZN(n18) );
  INV_X1 U63 ( .A(data_in[16]), .ZN(n59) );
  OAI22_X1 U64 ( .A1(n45), .A2(n58), .B1(net108243), .B2(n39), .ZN(n17) );
  INV_X1 U65 ( .A(data_in[17]), .ZN(n58) );
  OAI22_X1 U66 ( .A1(n46), .A2(n57), .B1(net108244), .B2(n39), .ZN(n16) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n57) );
  OAI22_X1 U68 ( .A1(n46), .A2(n56), .B1(net108245), .B2(n39), .ZN(n15) );
  INV_X1 U69 ( .A(data_in[19]), .ZN(n56) );
  OAI22_X1 U70 ( .A1(n46), .A2(n55), .B1(n37), .B2(n39), .ZN(n14) );
  INV_X1 U71 ( .A(data_in[20]), .ZN(n55) );
  OAI22_X1 U72 ( .A1(n46), .A2(n54), .B1(net108247), .B2(n39), .ZN(n13) );
  INV_X1 U73 ( .A(data_in[21]), .ZN(n54) );
  OAI22_X1 U74 ( .A1(n46), .A2(n53), .B1(net108248), .B2(n39), .ZN(n12) );
  INV_X1 U75 ( .A(data_in[22]), .ZN(n53) );
  OAI22_X1 U76 ( .A1(n47), .A2(n52), .B1(net108249), .B2(n39), .ZN(n11) );
  INV_X1 U77 ( .A(data_in[23]), .ZN(n52) );
  OAI22_X1 U78 ( .A1(n47), .A2(n51), .B1(net108250), .B2(n39), .ZN(n10) );
  INV_X1 U79 ( .A(data_in[24]), .ZN(n51) );
  OAI22_X1 U80 ( .A1(n45), .A2(n61), .B1(net108257), .B2(n39), .ZN(n2) );
  INV_X1 U81 ( .A(data_in[31]), .ZN(n61) );
  NAND2_X1 U82 ( .A1(load), .A2(enable), .ZN(n98) );
  INV_X1 U83 ( .A(reset), .ZN(n3) );
endmodule


module NRegister_N32_109 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n46), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n44), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n44), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n44), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n44), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n44), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n44), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n46), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n44), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n45), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n45), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n45), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n45), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n45), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n45), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n45), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n44), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n46), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n44), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n44), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n44), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n44), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n45), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n45), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n46), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n46), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n46), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n46), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n46), .Q(data_out[0]), 
        .QN(net108226) );
  INV_X1 U3 ( .A(n43), .ZN(n36) );
  INV_X1 U4 ( .A(n43), .ZN(n35) );
  BUF_X1 U5 ( .A(n92), .Z(n39) );
  BUF_X1 U6 ( .A(n92), .Z(n40) );
  BUF_X1 U7 ( .A(n92), .Z(n42) );
  BUF_X1 U8 ( .A(n92), .Z(n37) );
  BUF_X1 U9 ( .A(n92), .Z(n38) );
  BUF_X1 U10 ( .A(n92), .Z(n41) );
  BUF_X1 U11 ( .A(n92), .Z(n43) );
  BUF_X1 U12 ( .A(n47), .Z(n45) );
  BUF_X1 U13 ( .A(n47), .Z(n44) );
  BUF_X1 U14 ( .A(n47), .Z(n46) );
  OAI22_X1 U15 ( .A1(n38), .A2(n85), .B1(net108226), .B2(n36), .ZN(n34) );
  INV_X1 U16 ( .A(data_in[0]), .ZN(n85) );
  OAI22_X1 U17 ( .A1(n38), .A2(n84), .B1(net108227), .B2(n35), .ZN(n33) );
  INV_X1 U18 ( .A(data_in[1]), .ZN(n84) );
  OAI22_X1 U19 ( .A1(n37), .A2(n91), .B1(net108251), .B2(n36), .ZN(n9) );
  INV_X1 U20 ( .A(data_in[25]), .ZN(n91) );
  OAI22_X1 U21 ( .A1(n37), .A2(n90), .B1(net108252), .B2(n35), .ZN(n8) );
  INV_X1 U22 ( .A(data_in[26]), .ZN(n90) );
  OAI22_X1 U23 ( .A1(n37), .A2(n89), .B1(net108253), .B2(n36), .ZN(n7) );
  INV_X1 U24 ( .A(data_in[27]), .ZN(n89) );
  OAI22_X1 U25 ( .A1(n37), .A2(n88), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U26 ( .A(data_in[28]), .ZN(n88) );
  OAI22_X1 U27 ( .A1(n37), .A2(n87), .B1(net108255), .B2(n36), .ZN(n5) );
  INV_X1 U28 ( .A(data_in[29]), .ZN(n87) );
  OAI22_X1 U29 ( .A1(n38), .A2(n86), .B1(net108256), .B2(n35), .ZN(n4) );
  INV_X1 U30 ( .A(data_in[30]), .ZN(n86) );
  OAI22_X1 U31 ( .A1(n38), .A2(n83), .B1(net108228), .B2(n36), .ZN(n32) );
  INV_X1 U32 ( .A(data_in[2]), .ZN(n83) );
  OAI22_X1 U33 ( .A1(n38), .A2(n82), .B1(net108229), .B2(n36), .ZN(n31) );
  INV_X1 U34 ( .A(data_in[3]), .ZN(n82) );
  OAI22_X1 U35 ( .A1(n39), .A2(n81), .B1(net108230), .B2(n36), .ZN(n30) );
  INV_X1 U36 ( .A(data_in[4]), .ZN(n81) );
  OAI22_X1 U37 ( .A1(n39), .A2(n70), .B1(net108231), .B2(n36), .ZN(n29) );
  INV_X1 U38 ( .A(data_in[5]), .ZN(n70) );
  OAI22_X1 U39 ( .A1(n39), .A2(n67), .B1(net108232), .B2(n36), .ZN(n28) );
  INV_X1 U40 ( .A(data_in[6]), .ZN(n67) );
  OAI22_X1 U41 ( .A1(n39), .A2(n66), .B1(net108233), .B2(n36), .ZN(n27) );
  INV_X1 U42 ( .A(data_in[7]), .ZN(n66) );
  OAI22_X1 U43 ( .A1(n39), .A2(n65), .B1(net108234), .B2(n36), .ZN(n26) );
  INV_X1 U44 ( .A(data_in[8]), .ZN(n65) );
  OAI22_X1 U45 ( .A1(n40), .A2(n64), .B1(net108235), .B2(n36), .ZN(n25) );
  INV_X1 U46 ( .A(data_in[9]), .ZN(n64) );
  OAI22_X1 U47 ( .A1(n40), .A2(n63), .B1(net108236), .B2(n36), .ZN(n24) );
  INV_X1 U48 ( .A(data_in[10]), .ZN(n63) );
  OAI22_X1 U49 ( .A1(n40), .A2(n62), .B1(net108237), .B2(n36), .ZN(n23) );
  INV_X1 U50 ( .A(data_in[11]), .ZN(n62) );
  OAI22_X1 U51 ( .A1(n40), .A2(n61), .B1(net108238), .B2(n36), .ZN(n22) );
  INV_X1 U52 ( .A(data_in[12]), .ZN(n61) );
  OAI22_X1 U53 ( .A1(n40), .A2(n60), .B1(net108239), .B2(n36), .ZN(n21) );
  INV_X1 U54 ( .A(data_in[13]), .ZN(n60) );
  OAI22_X1 U55 ( .A1(n41), .A2(n59), .B1(net108240), .B2(n35), .ZN(n20) );
  INV_X1 U56 ( .A(data_in[14]), .ZN(n59) );
  OAI22_X1 U57 ( .A1(n41), .A2(n57), .B1(net108241), .B2(n35), .ZN(n19) );
  INV_X1 U58 ( .A(data_in[15]), .ZN(n57) );
  OAI22_X1 U59 ( .A1(n41), .A2(n56), .B1(net108242), .B2(n35), .ZN(n18) );
  INV_X1 U60 ( .A(data_in[16]), .ZN(n56) );
  OAI22_X1 U61 ( .A1(n41), .A2(n55), .B1(net108243), .B2(n35), .ZN(n17) );
  INV_X1 U62 ( .A(data_in[17]), .ZN(n55) );
  OAI22_X1 U63 ( .A1(n42), .A2(n54), .B1(net108244), .B2(n35), .ZN(n16) );
  INV_X1 U64 ( .A(data_in[18]), .ZN(n54) );
  OAI22_X1 U65 ( .A1(n42), .A2(n53), .B1(net108245), .B2(n35), .ZN(n15) );
  INV_X1 U66 ( .A(data_in[19]), .ZN(n53) );
  OAI22_X1 U67 ( .A1(n42), .A2(n52), .B1(net108246), .B2(n35), .ZN(n14) );
  INV_X1 U68 ( .A(data_in[20]), .ZN(n52) );
  OAI22_X1 U69 ( .A1(n42), .A2(n51), .B1(net108247), .B2(n35), .ZN(n13) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n51) );
  OAI22_X1 U71 ( .A1(n42), .A2(n50), .B1(net108248), .B2(n35), .ZN(n12) );
  INV_X1 U72 ( .A(data_in[22]), .ZN(n50) );
  OAI22_X1 U73 ( .A1(n43), .A2(n49), .B1(net108249), .B2(n35), .ZN(n11) );
  INV_X1 U74 ( .A(data_in[23]), .ZN(n49) );
  OAI22_X1 U75 ( .A1(n43), .A2(n48), .B1(net108250), .B2(n35), .ZN(n10) );
  INV_X1 U76 ( .A(data_in[24]), .ZN(n48) );
  OAI22_X1 U77 ( .A1(n41), .A2(n58), .B1(net108257), .B2(n35), .ZN(n2) );
  INV_X1 U78 ( .A(data_in[31]), .ZN(n58) );
  NAND2_X1 U79 ( .A1(load), .A2(enable), .ZN(n92) );
  INV_X1 U80 ( .A(reset), .ZN(n47) );
endmodule


module NRegister_N32_108 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n46), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n44), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n44), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n44), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n44), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n44), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n44), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n46), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n44), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n45), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n45), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n45), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n45), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n45), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n45), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n45), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n44), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n46), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n44), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n44), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n44), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n44), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n45), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n45), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n46), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n46), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n46), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n46), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n46), .Q(data_out[0]), 
        .QN(net108226) );
  INV_X1 U3 ( .A(n43), .ZN(n35) );
  BUF_X1 U4 ( .A(n92), .Z(n39) );
  BUF_X1 U5 ( .A(n92), .Z(n40) );
  BUF_X1 U6 ( .A(n92), .Z(n42) );
  BUF_X1 U7 ( .A(n92), .Z(n37) );
  BUF_X1 U8 ( .A(n92), .Z(n38) );
  BUF_X1 U9 ( .A(n92), .Z(n41) );
  BUF_X1 U10 ( .A(n92), .Z(n43) );
  BUF_X1 U11 ( .A(n47), .Z(n45) );
  BUF_X1 U12 ( .A(n47), .Z(n44) );
  BUF_X1 U13 ( .A(n47), .Z(n46) );
  OAI22_X1 U14 ( .A1(n38), .A2(n86), .B1(net108256), .B2(n36), .ZN(n4) );
  INV_X1 U15 ( .A(data_in[30]), .ZN(n86) );
  OAI22_X1 U16 ( .A1(n37), .A2(n87), .B1(net108255), .B2(n36), .ZN(n5) );
  INV_X1 U17 ( .A(data_in[29]), .ZN(n87) );
  OAI22_X1 U18 ( .A1(n37), .A2(n88), .B1(net108254), .B2(n36), .ZN(n6) );
  INV_X1 U19 ( .A(data_in[28]), .ZN(n88) );
  OAI22_X1 U20 ( .A1(n41), .A2(n58), .B1(net108257), .B2(n35), .ZN(n2) );
  INV_X1 U21 ( .A(data_in[31]), .ZN(n58) );
  OAI22_X1 U22 ( .A1(n37), .A2(n89), .B1(net108253), .B2(n36), .ZN(n7) );
  INV_X1 U23 ( .A(data_in[27]), .ZN(n89) );
  OAI22_X1 U24 ( .A1(n37), .A2(n90), .B1(net108252), .B2(n36), .ZN(n8) );
  INV_X1 U25 ( .A(data_in[26]), .ZN(n90) );
  OAI22_X1 U26 ( .A1(n37), .A2(n91), .B1(net108251), .B2(n36), .ZN(n9) );
  INV_X1 U27 ( .A(data_in[25]), .ZN(n91) );
  OAI22_X1 U28 ( .A1(n43), .A2(n48), .B1(net108250), .B2(n35), .ZN(n10) );
  INV_X1 U29 ( .A(data_in[24]), .ZN(n48) );
  OAI22_X1 U30 ( .A1(n43), .A2(n49), .B1(net108249), .B2(n35), .ZN(n11) );
  INV_X1 U31 ( .A(data_in[23]), .ZN(n49) );
  OAI22_X1 U32 ( .A1(n42), .A2(n50), .B1(net108248), .B2(n35), .ZN(n12) );
  INV_X1 U33 ( .A(data_in[22]), .ZN(n50) );
  OAI22_X1 U34 ( .A1(n42), .A2(n51), .B1(net108247), .B2(n35), .ZN(n13) );
  INV_X1 U35 ( .A(data_in[21]), .ZN(n51) );
  OAI22_X1 U36 ( .A1(n42), .A2(n52), .B1(net108246), .B2(n35), .ZN(n14) );
  INV_X1 U37 ( .A(data_in[20]), .ZN(n52) );
  OAI22_X1 U38 ( .A1(n41), .A2(n59), .B1(net108240), .B2(n35), .ZN(n20) );
  INV_X1 U39 ( .A(data_in[14]), .ZN(n59) );
  OAI22_X1 U40 ( .A1(n41), .A2(n57), .B1(net108241), .B2(n35), .ZN(n19) );
  INV_X1 U41 ( .A(data_in[15]), .ZN(n57) );
  OAI22_X1 U42 ( .A1(n41), .A2(n56), .B1(net108242), .B2(n35), .ZN(n18) );
  INV_X1 U43 ( .A(data_in[16]), .ZN(n56) );
  OAI22_X1 U44 ( .A1(n42), .A2(n53), .B1(net108245), .B2(n35), .ZN(n15) );
  INV_X1 U45 ( .A(data_in[19]), .ZN(n53) );
  OAI22_X1 U46 ( .A1(n42), .A2(n54), .B1(net108244), .B2(n35), .ZN(n16) );
  INV_X1 U47 ( .A(data_in[18]), .ZN(n54) );
  OAI22_X1 U48 ( .A1(n41), .A2(n55), .B1(net108243), .B2(n35), .ZN(n17) );
  INV_X1 U49 ( .A(data_in[17]), .ZN(n55) );
  OAI22_X1 U50 ( .A1(n39), .A2(n67), .B1(net108232), .B2(n35), .ZN(n28) );
  INV_X1 U51 ( .A(data_in[6]), .ZN(n67) );
  OAI22_X1 U52 ( .A1(n39), .A2(n66), .B1(net108233), .B2(n36), .ZN(n27) );
  INV_X1 U53 ( .A(data_in[7]), .ZN(n66) );
  OAI22_X1 U54 ( .A1(n39), .A2(n65), .B1(net108234), .B2(n35), .ZN(n26) );
  INV_X1 U55 ( .A(data_in[8]), .ZN(n65) );
  OAI22_X1 U56 ( .A1(n40), .A2(n64), .B1(net108235), .B2(n36), .ZN(n25) );
  INV_X1 U57 ( .A(data_in[9]), .ZN(n64) );
  OAI22_X1 U58 ( .A1(n40), .A2(n63), .B1(net108236), .B2(n35), .ZN(n24) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n63) );
  OAI22_X1 U60 ( .A1(n40), .A2(n62), .B1(net108237), .B2(n36), .ZN(n23) );
  INV_X1 U61 ( .A(data_in[11]), .ZN(n62) );
  OAI22_X1 U62 ( .A1(n40), .A2(n61), .B1(net108238), .B2(n35), .ZN(n22) );
  INV_X1 U63 ( .A(data_in[12]), .ZN(n61) );
  OAI22_X1 U64 ( .A1(n40), .A2(n60), .B1(net108239), .B2(n36), .ZN(n21) );
  INV_X1 U65 ( .A(data_in[13]), .ZN(n60) );
  OAI22_X1 U66 ( .A1(n38), .A2(n84), .B1(net108227), .B2(n36), .ZN(n33) );
  INV_X1 U67 ( .A(data_in[1]), .ZN(n84) );
  OAI22_X1 U68 ( .A1(n38), .A2(n83), .B1(net108228), .B2(n36), .ZN(n32) );
  INV_X1 U69 ( .A(data_in[2]), .ZN(n83) );
  OAI22_X1 U70 ( .A1(n38), .A2(n82), .B1(net108229), .B2(n36), .ZN(n31) );
  INV_X1 U71 ( .A(data_in[3]), .ZN(n82) );
  OAI22_X1 U72 ( .A1(n39), .A2(n81), .B1(net108230), .B2(n36), .ZN(n30) );
  INV_X1 U73 ( .A(data_in[4]), .ZN(n81) );
  OAI22_X1 U74 ( .A1(n39), .A2(n70), .B1(net108231), .B2(n36), .ZN(n29) );
  INV_X1 U75 ( .A(data_in[5]), .ZN(n70) );
  OAI22_X1 U76 ( .A1(n38), .A2(n85), .B1(net108226), .B2(n36), .ZN(n34) );
  INV_X1 U77 ( .A(data_in[0]), .ZN(n85) );
  NAND2_X1 U78 ( .A1(load), .A2(enable), .ZN(n92) );
  INV_X1 U79 ( .A(reset), .ZN(n47) );
  INV_X1 U80 ( .A(n43), .ZN(n36) );
endmodule


module NRegister_N32_107 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_106 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_105 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_104 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_103 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_102 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_101 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_100 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_99 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_98 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_97 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_96 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_95 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_94 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_93 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_92 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_91 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_90 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_89 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_88 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_87 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_86 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_85 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_84 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_83 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_82 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_81 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_80 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_79 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_78 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_77 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_76 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n80) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U17 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U18 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U22 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U23 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U24 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U25 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U26 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U27 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U28 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U29 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U30 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U31 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U32 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U33 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U34 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U35 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U36 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U37 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U38 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U39 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U40 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U41 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U42 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U44 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U45 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U46 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U47 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  NAND2_X1 U48 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_75 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_74 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_73 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_72 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_71 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_70 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_69 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_68 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_67 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_66 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_65 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_64 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_63 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_62 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_61 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_60 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_59 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_58 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_57 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_56 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_55 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_54 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_53 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_52 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_51 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_50 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_49 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_48 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_47 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_46 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_45 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_44 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n80) );
  BUF_X1 U8 ( .A(n81), .Z(n39) );
  BUF_X1 U9 ( .A(n81), .Z(n40) );
  BUF_X1 U10 ( .A(n81), .Z(n42) );
  BUF_X1 U11 ( .A(n81), .Z(n37) );
  BUF_X1 U12 ( .A(n81), .Z(n38) );
  BUF_X1 U13 ( .A(n81), .Z(n41) );
  BUF_X1 U14 ( .A(n81), .Z(n43) );
  OAI22_X1 U15 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  OAI22_X1 U16 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  OAI22_X1 U18 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U21 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U22 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U23 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U24 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U25 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U26 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U27 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U28 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U29 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n35), .ZN(n21) );
  OAI22_X1 U30 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U31 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U32 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U34 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U35 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n35), .ZN(n29) );
  OAI22_X1 U36 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U37 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n35), .ZN(n27) );
  OAI22_X1 U38 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U39 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n35), .ZN(n25) );
  OAI22_X1 U40 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U41 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U42 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U43 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n36), .ZN(n33) );
  OAI22_X1 U44 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U45 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U46 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  NAND2_X1 U47 ( .A1(load), .A2(enable), .ZN(n81) );
  INV_X1 U48 ( .A(n43), .ZN(n36) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_41 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, net108226, net108227, net108228, net108229,
         net108230, net108231, net108232, net108233, net108234, net108235,
         net108236, net108237, net108238, net108239, net108240, net108241,
         net108242, net108243, net108244, net108245, net108246, net108247,
         net108248, net108249, net108250, net108251, net108252, net108253,
         net108254, net108255, net108256, net108257, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n70, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n44), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n46), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n46), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n46), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n45), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n45), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n45), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n44), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n45), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n45), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n45), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n45), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n45), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n45), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n45), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n45), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n46), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n44), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n46), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n44), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n46), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n46), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n46), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n44), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n44), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n44), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n44), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n44), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n44), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n44), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n44), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n3), .Z(n45) );
  BUF_X1 U4 ( .A(n3), .Z(n44) );
  BUF_X1 U5 ( .A(n3), .Z(n46) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n3) );
  BUF_X1 U9 ( .A(n90), .Z(n39) );
  BUF_X1 U10 ( .A(n90), .Z(n40) );
  BUF_X1 U11 ( .A(n90), .Z(n42) );
  BUF_X1 U12 ( .A(n90), .Z(n37) );
  BUF_X1 U13 ( .A(n90), .Z(n38) );
  BUF_X1 U14 ( .A(n90), .Z(n41) );
  BUF_X1 U15 ( .A(n90), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n83), .B1(net108226), .B2(n36), .ZN(n34) );
  INV_X1 U17 ( .A(data_in[0]), .ZN(n83) );
  OAI22_X1 U18 ( .A1(n38), .A2(n82), .B1(net108227), .B2(n35), .ZN(n33) );
  INV_X1 U19 ( .A(data_in[1]), .ZN(n82) );
  OAI22_X1 U20 ( .A1(n37), .A2(n89), .B1(net108251), .B2(n36), .ZN(n9) );
  INV_X1 U21 ( .A(data_in[25]), .ZN(n89) );
  OAI22_X1 U22 ( .A1(n37), .A2(n88), .B1(net108252), .B2(n35), .ZN(n8) );
  INV_X1 U23 ( .A(data_in[26]), .ZN(n88) );
  OAI22_X1 U24 ( .A1(n37), .A2(n87), .B1(net108253), .B2(n36), .ZN(n7) );
  INV_X1 U25 ( .A(data_in[27]), .ZN(n87) );
  OAI22_X1 U26 ( .A1(n37), .A2(n86), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U27 ( .A(data_in[28]), .ZN(n86) );
  OAI22_X1 U28 ( .A1(n37), .A2(n85), .B1(net108255), .B2(n36), .ZN(n5) );
  INV_X1 U29 ( .A(data_in[29]), .ZN(n85) );
  OAI22_X1 U30 ( .A1(n38), .A2(n84), .B1(net108256), .B2(n35), .ZN(n4) );
  INV_X1 U31 ( .A(data_in[30]), .ZN(n84) );
  OAI22_X1 U32 ( .A1(n38), .A2(n81), .B1(net108228), .B2(n36), .ZN(n32) );
  INV_X1 U33 ( .A(data_in[2]), .ZN(n81) );
  OAI22_X1 U34 ( .A1(n38), .A2(n80), .B1(net108229), .B2(n36), .ZN(n31) );
  INV_X1 U35 ( .A(data_in[3]), .ZN(n80) );
  OAI22_X1 U36 ( .A1(n39), .A2(n70), .B1(net108230), .B2(n36), .ZN(n30) );
  INV_X1 U37 ( .A(data_in[4]), .ZN(n70) );
  OAI22_X1 U38 ( .A1(n39), .A2(n67), .B1(net108231), .B2(n36), .ZN(n29) );
  INV_X1 U39 ( .A(data_in[5]), .ZN(n67) );
  OAI22_X1 U40 ( .A1(n39), .A2(n66), .B1(net108232), .B2(n36), .ZN(n28) );
  INV_X1 U41 ( .A(data_in[6]), .ZN(n66) );
  OAI22_X1 U42 ( .A1(n39), .A2(n65), .B1(net108233), .B2(n36), .ZN(n27) );
  INV_X1 U43 ( .A(data_in[7]), .ZN(n65) );
  OAI22_X1 U44 ( .A1(n39), .A2(n64), .B1(net108234), .B2(n36), .ZN(n26) );
  INV_X1 U45 ( .A(data_in[8]), .ZN(n64) );
  OAI22_X1 U46 ( .A1(n40), .A2(n63), .B1(net108235), .B2(n36), .ZN(n25) );
  INV_X1 U47 ( .A(data_in[9]), .ZN(n63) );
  OAI22_X1 U48 ( .A1(n40), .A2(n62), .B1(net108236), .B2(n36), .ZN(n24) );
  INV_X1 U49 ( .A(data_in[10]), .ZN(n62) );
  OAI22_X1 U50 ( .A1(n40), .A2(n61), .B1(net108237), .B2(n36), .ZN(n23) );
  INV_X1 U51 ( .A(data_in[11]), .ZN(n61) );
  OAI22_X1 U52 ( .A1(n40), .A2(n60), .B1(net108238), .B2(n36), .ZN(n22) );
  INV_X1 U53 ( .A(data_in[12]), .ZN(n60) );
  OAI22_X1 U54 ( .A1(n40), .A2(n59), .B1(net108239), .B2(n36), .ZN(n21) );
  INV_X1 U55 ( .A(data_in[13]), .ZN(n59) );
  OAI22_X1 U56 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  INV_X1 U57 ( .A(data_in[14]), .ZN(n58) );
  OAI22_X1 U58 ( .A1(n41), .A2(n56), .B1(net108241), .B2(n35), .ZN(n19) );
  INV_X1 U59 ( .A(data_in[15]), .ZN(n56) );
  OAI22_X1 U60 ( .A1(n41), .A2(n55), .B1(net108242), .B2(n35), .ZN(n18) );
  INV_X1 U61 ( .A(data_in[16]), .ZN(n55) );
  OAI22_X1 U62 ( .A1(n41), .A2(n54), .B1(net108243), .B2(n35), .ZN(n17) );
  INV_X1 U63 ( .A(data_in[17]), .ZN(n54) );
  OAI22_X1 U64 ( .A1(n42), .A2(n53), .B1(net108244), .B2(n35), .ZN(n16) );
  INV_X1 U65 ( .A(data_in[18]), .ZN(n53) );
  OAI22_X1 U66 ( .A1(n42), .A2(n52), .B1(net108245), .B2(n35), .ZN(n15) );
  INV_X1 U67 ( .A(data_in[19]), .ZN(n52) );
  OAI22_X1 U68 ( .A1(n42), .A2(n51), .B1(net108246), .B2(n35), .ZN(n14) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n51) );
  OAI22_X1 U70 ( .A1(n42), .A2(n50), .B1(net108247), .B2(n35), .ZN(n13) );
  INV_X1 U71 ( .A(data_in[21]), .ZN(n50) );
  OAI22_X1 U72 ( .A1(n42), .A2(n49), .B1(net108248), .B2(n35), .ZN(n12) );
  INV_X1 U73 ( .A(data_in[22]), .ZN(n49) );
  OAI22_X1 U74 ( .A1(n43), .A2(n48), .B1(net108249), .B2(n35), .ZN(n11) );
  INV_X1 U75 ( .A(data_in[23]), .ZN(n48) );
  OAI22_X1 U76 ( .A1(n43), .A2(n47), .B1(net108250), .B2(n35), .ZN(n10) );
  INV_X1 U77 ( .A(data_in[24]), .ZN(n47) );
  OAI22_X1 U78 ( .A1(n41), .A2(n57), .B1(net108257), .B2(n35), .ZN(n2) );
  INV_X1 U79 ( .A(data_in[31]), .ZN(n57) );
  NAND2_X1 U80 ( .A1(load), .A2(enable), .ZN(n90) );
endmodule


module NRegister_N32_34 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, net108226, net108227, net108228, net108229,
         net108230, net108231, net108232, net108233, net108234, net108235,
         net108236, net108237, net108238, net108239, net108240, net108241,
         net108242, net108243, net108244, net108245, net108246, net108247,
         net108248, net108249, net108250, net108251, net108252, net108253,
         net108254, net108255, net108256, net108257, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n70, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n44), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n46), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n46), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n46), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n45), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n45), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n45), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n44), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n45), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n45), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n45), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n45), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n45), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n45), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n45), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n45), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n46), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n44), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n46), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n44), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n46), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n46), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n46), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n44), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n44), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n44), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n44), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n44), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n44), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n44), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n44), .Q(data_out[0]), 
        .QN(net108226) );
  INV_X1 U3 ( .A(n43), .ZN(n35) );
  BUF_X1 U4 ( .A(n90), .Z(n39) );
  BUF_X1 U5 ( .A(n90), .Z(n40) );
  BUF_X1 U6 ( .A(n90), .Z(n42) );
  BUF_X1 U7 ( .A(n90), .Z(n37) );
  BUF_X1 U8 ( .A(n90), .Z(n38) );
  BUF_X1 U9 ( .A(n90), .Z(n41) );
  BUF_X1 U10 ( .A(n90), .Z(n43) );
  BUF_X1 U11 ( .A(n3), .Z(n45) );
  BUF_X1 U12 ( .A(n3), .Z(n44) );
  BUF_X1 U13 ( .A(n3), .Z(n46) );
  OAI22_X1 U14 ( .A1(n38), .A2(n83), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U15 ( .A1(n38), .A2(n81), .B1(net108228), .B2(n35), .ZN(n32) );
  INV_X1 U16 ( .A(data_in[2]), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n40), .A2(n60), .B1(net108238), .B2(n35), .ZN(n22) );
  INV_X1 U18 ( .A(data_in[12]), .ZN(n60) );
  OAI22_X1 U19 ( .A1(n40), .A2(n59), .B1(net108239), .B2(n35), .ZN(n21) );
  INV_X1 U20 ( .A(data_in[13]), .ZN(n59) );
  OAI22_X1 U21 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  INV_X1 U22 ( .A(data_in[14]), .ZN(n58) );
  OAI22_X1 U23 ( .A1(n41), .A2(n54), .B1(net108243), .B2(n36), .ZN(n17) );
  INV_X1 U24 ( .A(data_in[17]), .ZN(n54) );
  OAI22_X1 U25 ( .A1(n41), .A2(n57), .B1(net108257), .B2(n35), .ZN(n2) );
  INV_X1 U26 ( .A(data_in[31]), .ZN(n57) );
  OAI22_X1 U27 ( .A1(n39), .A2(n66), .B1(net108232), .B2(n35), .ZN(n28) );
  INV_X1 U28 ( .A(data_in[6]), .ZN(n66) );
  OAI22_X1 U29 ( .A1(n39), .A2(n70), .B1(net108230), .B2(n35), .ZN(n30) );
  INV_X1 U30 ( .A(data_in[4]), .ZN(n70) );
  OAI22_X1 U31 ( .A1(n38), .A2(n84), .B1(net108256), .B2(n36), .ZN(n4) );
  INV_X1 U32 ( .A(data_in[30]), .ZN(n84) );
  OAI22_X1 U33 ( .A1(n42), .A2(n51), .B1(net108246), .B2(n36), .ZN(n14) );
  INV_X1 U34 ( .A(data_in[20]), .ZN(n51) );
  OAI22_X1 U35 ( .A1(n37), .A2(n86), .B1(net108254), .B2(n36), .ZN(n6) );
  INV_X1 U36 ( .A(data_in[28]), .ZN(n86) );
  OAI22_X1 U37 ( .A1(n39), .A2(n64), .B1(net108234), .B2(n35), .ZN(n26) );
  INV_X1 U38 ( .A(data_in[8]), .ZN(n64) );
  OAI22_X1 U39 ( .A1(n42), .A2(n49), .B1(net108248), .B2(n35), .ZN(n12) );
  INV_X1 U40 ( .A(data_in[22]), .ZN(n49) );
  OAI22_X1 U41 ( .A1(n37), .A2(n88), .B1(net108252), .B2(n36), .ZN(n8) );
  INV_X1 U42 ( .A(data_in[26]), .ZN(n88) );
  OAI22_X1 U43 ( .A1(n41), .A2(n55), .B1(net108242), .B2(n36), .ZN(n18) );
  INV_X1 U44 ( .A(data_in[16]), .ZN(n55) );
  OAI22_X1 U45 ( .A1(n38), .A2(n80), .B1(net108229), .B2(n35), .ZN(n31) );
  INV_X1 U46 ( .A(data_in[3]), .ZN(n80) );
  OAI22_X1 U47 ( .A1(n39), .A2(n65), .B1(net108233), .B2(n35), .ZN(n27) );
  INV_X1 U48 ( .A(data_in[7]), .ZN(n65) );
  OAI22_X1 U49 ( .A1(n39), .A2(n67), .B1(net108231), .B2(n35), .ZN(n29) );
  INV_X1 U50 ( .A(data_in[5]), .ZN(n67) );
  OAI22_X1 U51 ( .A1(n42), .A2(n50), .B1(net108247), .B2(n35), .ZN(n13) );
  INV_X1 U52 ( .A(data_in[21]), .ZN(n50) );
  OAI22_X1 U53 ( .A1(n37), .A2(n85), .B1(net108255), .B2(n36), .ZN(n5) );
  INV_X1 U54 ( .A(data_in[29]), .ZN(n85) );
  OAI22_X1 U55 ( .A1(n41), .A2(n56), .B1(net108241), .B2(n36), .ZN(n19) );
  INV_X1 U56 ( .A(data_in[15]), .ZN(n56) );
  OAI22_X1 U57 ( .A1(n40), .A2(n63), .B1(net108235), .B2(n35), .ZN(n25) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n63) );
  OAI22_X1 U59 ( .A1(n43), .A2(n48), .B1(net108249), .B2(n36), .ZN(n11) );
  INV_X1 U60 ( .A(data_in[23]), .ZN(n48) );
  OAI22_X1 U61 ( .A1(n37), .A2(n87), .B1(net108253), .B2(n36), .ZN(n7) );
  INV_X1 U62 ( .A(data_in[27]), .ZN(n87) );
  OAI22_X1 U63 ( .A1(n40), .A2(n62), .B1(net108236), .B2(n35), .ZN(n24) );
  INV_X1 U64 ( .A(data_in[10]), .ZN(n62) );
  OAI22_X1 U65 ( .A1(n43), .A2(n47), .B1(net108250), .B2(n36), .ZN(n10) );
  INV_X1 U66 ( .A(data_in[24]), .ZN(n47) );
  OAI22_X1 U67 ( .A1(n42), .A2(n53), .B1(net108244), .B2(n36), .ZN(n16) );
  INV_X1 U68 ( .A(data_in[18]), .ZN(n53) );
  OAI22_X1 U69 ( .A1(n37), .A2(n89), .B1(net108251), .B2(n36), .ZN(n9) );
  INV_X1 U70 ( .A(data_in[25]), .ZN(n89) );
  OAI22_X1 U71 ( .A1(n40), .A2(n61), .B1(net108237), .B2(n35), .ZN(n23) );
  INV_X1 U72 ( .A(data_in[11]), .ZN(n61) );
  OAI22_X1 U73 ( .A1(n42), .A2(n52), .B1(net108245), .B2(n36), .ZN(n15) );
  INV_X1 U74 ( .A(data_in[19]), .ZN(n52) );
  OAI22_X1 U75 ( .A1(n38), .A2(n82), .B1(net108227), .B2(n36), .ZN(n33) );
  INV_X1 U76 ( .A(data_in[1]), .ZN(n82) );
  NAND2_X1 U77 ( .A1(load), .A2(enable), .ZN(n90) );
  INV_X1 U78 ( .A(reset), .ZN(n3) );
  INV_X1 U79 ( .A(data_in[0]), .ZN(n83) );
  INV_X1 U80 ( .A(n43), .ZN(n36) );
endmodule


module NRegister_N32_30 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_29 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_28 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_27 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_26 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_25 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_23 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_22 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_21 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_20 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_19 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_18 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_17 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_16 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_15 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_13 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_12 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_11 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_10 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_9 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_8 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_7 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_6 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_4 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  OAI22_X1 U20 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n35), .ZN(n7) );
  OAI22_X1 U21 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U22 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U23 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U24 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U25 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U26 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U27 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U28 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U29 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U30 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U31 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  OAI22_X1 U32 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U33 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U34 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U35 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U36 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U37 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U38 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U39 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U40 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U41 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U42 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U43 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U44 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U45 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U48 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_3 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U20 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U21 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U22 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U23 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U24 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U25 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U26 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U27 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U28 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U29 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U30 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U31 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U32 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U33 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U34 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U35 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U36 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U37 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U38 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U39 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U40 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U41 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U42 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U43 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U44 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U45 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U48 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_2 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U20 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U21 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U22 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U23 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U24 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U25 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U26 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U27 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U28 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U29 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U30 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U31 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U32 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U33 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U34 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U35 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U36 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U37 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U38 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U39 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U40 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U41 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U42 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U43 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U44 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U45 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U48 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_1 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n77), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n77), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n77), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n79), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n77), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n78), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n78), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n78), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n78), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n78), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n78), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n78), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n79), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n77), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n77), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n77), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n77), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n79), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n79), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108226), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108227), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n70), .B1(net108251), .B2(n36), .ZN(n9) );
  OAI22_X1 U20 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n35), .ZN(n8) );
  OAI22_X1 U21 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  OAI22_X1 U22 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n35), .ZN(n6) );
  OAI22_X1 U23 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  OAI22_X1 U24 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n35), .ZN(n4) );
  OAI22_X1 U25 ( .A1(n38), .A2(n46), .B1(net108228), .B2(n36), .ZN(n32) );
  OAI22_X1 U26 ( .A1(n38), .A2(n47), .B1(net108229), .B2(n36), .ZN(n31) );
  OAI22_X1 U27 ( .A1(n39), .A2(n48), .B1(net108230), .B2(n36), .ZN(n30) );
  OAI22_X1 U28 ( .A1(n39), .A2(n49), .B1(net108231), .B2(n36), .ZN(n29) );
  OAI22_X1 U29 ( .A1(n39), .A2(n50), .B1(net108232), .B2(n36), .ZN(n28) );
  OAI22_X1 U30 ( .A1(n39), .A2(n51), .B1(net108233), .B2(n36), .ZN(n27) );
  OAI22_X1 U31 ( .A1(n39), .A2(n52), .B1(net108234), .B2(n36), .ZN(n26) );
  OAI22_X1 U32 ( .A1(n40), .A2(n53), .B1(net108235), .B2(n36), .ZN(n25) );
  OAI22_X1 U33 ( .A1(n40), .A2(n54), .B1(net108236), .B2(n36), .ZN(n24) );
  OAI22_X1 U34 ( .A1(n40), .A2(n55), .B1(net108237), .B2(n36), .ZN(n23) );
  OAI22_X1 U35 ( .A1(n40), .A2(n56), .B1(net108238), .B2(n36), .ZN(n22) );
  OAI22_X1 U36 ( .A1(n40), .A2(n57), .B1(net108239), .B2(n36), .ZN(n21) );
  OAI22_X1 U37 ( .A1(n41), .A2(n58), .B1(net108240), .B2(n35), .ZN(n20) );
  OAI22_X1 U38 ( .A1(n41), .A2(n59), .B1(net108241), .B2(n35), .ZN(n19) );
  OAI22_X1 U39 ( .A1(n41), .A2(n60), .B1(net108242), .B2(n35), .ZN(n18) );
  OAI22_X1 U40 ( .A1(n41), .A2(n61), .B1(net108243), .B2(n35), .ZN(n17) );
  OAI22_X1 U41 ( .A1(n42), .A2(n62), .B1(net108244), .B2(n35), .ZN(n16) );
  OAI22_X1 U42 ( .A1(n42), .A2(n63), .B1(net108245), .B2(n35), .ZN(n15) );
  OAI22_X1 U43 ( .A1(n42), .A2(n64), .B1(net108246), .B2(n35), .ZN(n14) );
  OAI22_X1 U44 ( .A1(n42), .A2(n65), .B1(net108247), .B2(n35), .ZN(n13) );
  OAI22_X1 U45 ( .A1(n42), .A2(n66), .B1(net108248), .B2(n35), .ZN(n12) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108249), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n43), .A2(n69), .B1(net108250), .B2(n35), .ZN(n10) );
  OAI22_X1 U48 ( .A1(n41), .A2(n76), .B1(net108257), .B2(n35), .ZN(n2) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_116 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108194, net108195, net108196, net108197, net108198,
         net108199, net108200, net108201, net108202, net108203, net108204,
         net108205, net108206, net108207, net108208, net108209, net108210,
         net108211, net108212, net108213, net108214, net108215, net108216,
         net108217, net108218, net108219, net108220, net108221, net108222,
         net108223, net108224, net108225, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n46), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n46), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n46), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n44), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n46), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n44), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n44), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n44), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n46), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n44), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n44), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n44), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n44), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n44), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n44), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n44), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n44), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n45), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n45), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n45), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n45), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n45), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n45), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n45), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n45), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n45), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n46), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n46), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n46), .Q(data_out[0]), 
        .QN(net108194) );
  BUF_X1 U3 ( .A(n47), .Z(n45) );
  BUF_X1 U4 ( .A(n47), .Z(n44) );
  BUF_X1 U5 ( .A(n47), .Z(n46) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n47) );
  BUF_X1 U9 ( .A(n92), .Z(n39) );
  BUF_X1 U10 ( .A(n92), .Z(n40) );
  BUF_X1 U11 ( .A(n92), .Z(n42) );
  BUF_X1 U12 ( .A(n92), .Z(n37) );
  BUF_X1 U13 ( .A(n92), .Z(n38) );
  BUF_X1 U14 ( .A(n92), .Z(n41) );
  BUF_X1 U15 ( .A(n92), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n85), .B1(net108194), .B2(n36), .ZN(n34) );
  INV_X1 U17 ( .A(data_in[0]), .ZN(n85) );
  OAI22_X1 U18 ( .A1(n38), .A2(n84), .B1(net108195), .B2(n35), .ZN(n33) );
  INV_X1 U19 ( .A(data_in[1]), .ZN(n84) );
  OAI22_X1 U20 ( .A1(n37), .A2(n91), .B1(net108219), .B2(n36), .ZN(n9) );
  INV_X1 U21 ( .A(data_in[25]), .ZN(n91) );
  OAI22_X1 U22 ( .A1(n37), .A2(n90), .B1(net108220), .B2(n35), .ZN(n8) );
  INV_X1 U23 ( .A(data_in[26]), .ZN(n90) );
  OAI22_X1 U24 ( .A1(n37), .A2(n89), .B1(net108221), .B2(n36), .ZN(n7) );
  INV_X1 U25 ( .A(data_in[27]), .ZN(n89) );
  OAI22_X1 U26 ( .A1(n37), .A2(n88), .B1(net108222), .B2(n35), .ZN(n6) );
  INV_X1 U27 ( .A(data_in[28]), .ZN(n88) );
  OAI22_X1 U28 ( .A1(n37), .A2(n87), .B1(net108223), .B2(n36), .ZN(n5) );
  INV_X1 U29 ( .A(data_in[29]), .ZN(n87) );
  OAI22_X1 U30 ( .A1(n38), .A2(n86), .B1(net108224), .B2(n35), .ZN(n4) );
  INV_X1 U31 ( .A(data_in[30]), .ZN(n86) );
  OAI22_X1 U32 ( .A1(n38), .A2(n83), .B1(net108196), .B2(n36), .ZN(n32) );
  INV_X1 U33 ( .A(data_in[2]), .ZN(n83) );
  OAI22_X1 U34 ( .A1(n38), .A2(n82), .B1(net108197), .B2(n36), .ZN(n31) );
  INV_X1 U35 ( .A(data_in[3]), .ZN(n82) );
  OAI22_X1 U36 ( .A1(n39), .A2(n81), .B1(net108198), .B2(n36), .ZN(n30) );
  INV_X1 U37 ( .A(data_in[4]), .ZN(n81) );
  OAI22_X1 U38 ( .A1(n39), .A2(n70), .B1(net108199), .B2(n36), .ZN(n29) );
  INV_X1 U39 ( .A(data_in[5]), .ZN(n70) );
  OAI22_X1 U40 ( .A1(n39), .A2(n67), .B1(net108200), .B2(n36), .ZN(n28) );
  INV_X1 U41 ( .A(data_in[6]), .ZN(n67) );
  OAI22_X1 U42 ( .A1(n39), .A2(n66), .B1(net108201), .B2(n36), .ZN(n27) );
  INV_X1 U43 ( .A(data_in[7]), .ZN(n66) );
  OAI22_X1 U44 ( .A1(n39), .A2(n65), .B1(net108202), .B2(n36), .ZN(n26) );
  INV_X1 U45 ( .A(data_in[8]), .ZN(n65) );
  OAI22_X1 U46 ( .A1(n40), .A2(n64), .B1(net108203), .B2(n36), .ZN(n25) );
  INV_X1 U47 ( .A(data_in[9]), .ZN(n64) );
  OAI22_X1 U48 ( .A1(n40), .A2(n63), .B1(net108204), .B2(n36), .ZN(n24) );
  INV_X1 U49 ( .A(data_in[10]), .ZN(n63) );
  OAI22_X1 U50 ( .A1(n40), .A2(n62), .B1(net108205), .B2(n36), .ZN(n23) );
  INV_X1 U51 ( .A(data_in[11]), .ZN(n62) );
  OAI22_X1 U52 ( .A1(n40), .A2(n61), .B1(net108206), .B2(n36), .ZN(n22) );
  INV_X1 U53 ( .A(data_in[12]), .ZN(n61) );
  OAI22_X1 U54 ( .A1(n40), .A2(n60), .B1(net108207), .B2(n36), .ZN(n21) );
  INV_X1 U55 ( .A(data_in[13]), .ZN(n60) );
  OAI22_X1 U56 ( .A1(n41), .A2(n59), .B1(net108208), .B2(n35), .ZN(n20) );
  INV_X1 U57 ( .A(data_in[14]), .ZN(n59) );
  OAI22_X1 U58 ( .A1(n41), .A2(n57), .B1(net108209), .B2(n35), .ZN(n19) );
  INV_X1 U59 ( .A(data_in[15]), .ZN(n57) );
  OAI22_X1 U60 ( .A1(n41), .A2(n56), .B1(net108210), .B2(n35), .ZN(n18) );
  INV_X1 U61 ( .A(data_in[16]), .ZN(n56) );
  OAI22_X1 U62 ( .A1(n41), .A2(n55), .B1(net108211), .B2(n35), .ZN(n17) );
  INV_X1 U63 ( .A(data_in[17]), .ZN(n55) );
  OAI22_X1 U64 ( .A1(n42), .A2(n54), .B1(net108212), .B2(n35), .ZN(n16) );
  INV_X1 U65 ( .A(data_in[18]), .ZN(n54) );
  OAI22_X1 U66 ( .A1(n42), .A2(n53), .B1(net108213), .B2(n35), .ZN(n15) );
  INV_X1 U67 ( .A(data_in[19]), .ZN(n53) );
  OAI22_X1 U68 ( .A1(n42), .A2(n52), .B1(net108214), .B2(n35), .ZN(n14) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n52) );
  OAI22_X1 U70 ( .A1(n42), .A2(n51), .B1(net108215), .B2(n35), .ZN(n13) );
  INV_X1 U71 ( .A(data_in[21]), .ZN(n51) );
  OAI22_X1 U72 ( .A1(n42), .A2(n50), .B1(net108216), .B2(n35), .ZN(n12) );
  INV_X1 U73 ( .A(data_in[22]), .ZN(n50) );
  OAI22_X1 U74 ( .A1(n43), .A2(n49), .B1(net108217), .B2(n35), .ZN(n11) );
  INV_X1 U75 ( .A(data_in[23]), .ZN(n49) );
  OAI22_X1 U76 ( .A1(n43), .A2(n48), .B1(net108218), .B2(n35), .ZN(n10) );
  INV_X1 U77 ( .A(data_in[24]), .ZN(n48) );
  OAI22_X1 U78 ( .A1(n41), .A2(n58), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U79 ( .A(data_in[31]), .ZN(n58) );
  NAND2_X1 U80 ( .A1(load), .A2(enable), .ZN(n92) );
endmodule


module NRegister_N32_114 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, net108194, net108195, net108196, net108197,
         net108198, net108199, net108200, net108201, net108202, net108203,
         net108204, net108205, net108206, net108207, net108208, net108209,
         net108210, net108211, net108212, net108213, net108214, net108215,
         net108216, net108217, net108218, net108219, net108220, net108221,
         net108222, net108223, net108224, net108225, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n70, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n44), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n44), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n44), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n46), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n44), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n46), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n46), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n46), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n44), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n46), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n46), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n46), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n45), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n45), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n45), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n45), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n45), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n44), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n44), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n44), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n44), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n44), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n44), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n44), .Q(data_out[0]), 
        .QN(net108194) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n45), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n45), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n46), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n45), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n45), .Q(data_out[18]), 
        .QN(net108212) );
  INV_X1 U3 ( .A(n43), .ZN(n35) );
  INV_X1 U4 ( .A(n43), .ZN(n36) );
  BUF_X1 U5 ( .A(n90), .Z(n39) );
  BUF_X1 U6 ( .A(n90), .Z(n42) );
  BUF_X1 U7 ( .A(n90), .Z(n37) );
  BUF_X1 U8 ( .A(n90), .Z(n38) );
  BUF_X1 U9 ( .A(n90), .Z(n41) );
  BUF_X1 U10 ( .A(n90), .Z(n43) );
  BUF_X1 U11 ( .A(n90), .Z(n40) );
  BUF_X1 U12 ( .A(n3), .Z(n45) );
  BUF_X1 U13 ( .A(n3), .Z(n44) );
  BUF_X1 U14 ( .A(n3), .Z(n46) );
  INV_X1 U15 ( .A(data_in[13]), .ZN(n59) );
  OAI22_X1 U16 ( .A1(n38), .A2(n83), .B1(net108194), .B2(n35), .ZN(n34) );
  INV_X1 U17 ( .A(data_in[0]), .ZN(n83) );
  OAI22_X1 U18 ( .A1(n38), .A2(n82), .B1(net108195), .B2(n36), .ZN(n33) );
  INV_X1 U19 ( .A(data_in[1]), .ZN(n82) );
  OAI22_X1 U20 ( .A1(n37), .A2(n89), .B1(net108219), .B2(n35), .ZN(n9) );
  INV_X1 U21 ( .A(data_in[25]), .ZN(n89) );
  OAI22_X1 U22 ( .A1(n37), .A2(n88), .B1(net108220), .B2(n36), .ZN(n8) );
  INV_X1 U23 ( .A(data_in[26]), .ZN(n88) );
  OAI22_X1 U24 ( .A1(n37), .A2(n87), .B1(net108221), .B2(n35), .ZN(n7) );
  INV_X1 U25 ( .A(data_in[27]), .ZN(n87) );
  OAI22_X1 U26 ( .A1(n37), .A2(n86), .B1(net108222), .B2(n36), .ZN(n6) );
  INV_X1 U27 ( .A(data_in[28]), .ZN(n86) );
  OAI22_X1 U28 ( .A1(n37), .A2(n85), .B1(net108223), .B2(n35), .ZN(n5) );
  INV_X1 U29 ( .A(data_in[29]), .ZN(n85) );
  OAI22_X1 U30 ( .A1(n38), .A2(n84), .B1(net108224), .B2(n36), .ZN(n4) );
  INV_X1 U31 ( .A(data_in[30]), .ZN(n84) );
  OAI22_X1 U32 ( .A1(n41), .A2(n55), .B1(net108210), .B2(n35), .ZN(n18) );
  OAI22_X1 U33 ( .A1(n41), .A2(n58), .B1(net108208), .B2(n35), .ZN(n20) );
  INV_X1 U34 ( .A(data_in[14]), .ZN(n58) );
  OAI22_X1 U35 ( .A1(n41), .A2(n56), .B1(net108209), .B2(n35), .ZN(n19) );
  INV_X1 U36 ( .A(data_in[15]), .ZN(n56) );
  OAI22_X1 U37 ( .A1(n41), .A2(n54), .B1(net108211), .B2(n35), .ZN(n17) );
  OAI22_X1 U38 ( .A1(n42), .A2(n53), .B1(net108212), .B2(n35), .ZN(n16) );
  INV_X1 U39 ( .A(data_in[18]), .ZN(n53) );
  OAI22_X1 U40 ( .A1(n42), .A2(n52), .B1(net108213), .B2(n35), .ZN(n15) );
  INV_X1 U41 ( .A(data_in[19]), .ZN(n52) );
  OAI22_X1 U42 ( .A1(n42), .A2(n51), .B1(net108214), .B2(n35), .ZN(n14) );
  OAI22_X1 U43 ( .A1(n42), .A2(n50), .B1(net108215), .B2(n35), .ZN(n13) );
  INV_X1 U44 ( .A(data_in[21]), .ZN(n50) );
  OAI22_X1 U45 ( .A1(n42), .A2(n49), .B1(net108216), .B2(n35), .ZN(n12) );
  INV_X1 U46 ( .A(data_in[22]), .ZN(n49) );
  OAI22_X1 U47 ( .A1(n43), .A2(n48), .B1(net108217), .B2(n35), .ZN(n11) );
  INV_X1 U48 ( .A(data_in[23]), .ZN(n48) );
  OAI22_X1 U49 ( .A1(n43), .A2(n47), .B1(net108218), .B2(n35), .ZN(n10) );
  INV_X1 U50 ( .A(data_in[24]), .ZN(n47) );
  OAI22_X1 U51 ( .A1(n41), .A2(n57), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U52 ( .A(data_in[31]), .ZN(n57) );
  OAI22_X1 U53 ( .A1(n38), .A2(n81), .B1(net108196), .B2(n36), .ZN(n32) );
  INV_X1 U54 ( .A(data_in[2]), .ZN(n81) );
  OAI22_X1 U55 ( .A1(n38), .A2(n80), .B1(net108197), .B2(n36), .ZN(n31) );
  INV_X1 U56 ( .A(data_in[3]), .ZN(n80) );
  OAI22_X1 U57 ( .A1(n39), .A2(n70), .B1(net108198), .B2(n36), .ZN(n30) );
  INV_X1 U58 ( .A(data_in[4]), .ZN(n70) );
  OAI22_X1 U59 ( .A1(n39), .A2(n67), .B1(net108199), .B2(n36), .ZN(n29) );
  INV_X1 U60 ( .A(data_in[5]), .ZN(n67) );
  OAI22_X1 U61 ( .A1(n39), .A2(n66), .B1(net108200), .B2(n36), .ZN(n28) );
  INV_X1 U62 ( .A(data_in[6]), .ZN(n66) );
  OAI22_X1 U63 ( .A1(n39), .A2(n65), .B1(net108201), .B2(n36), .ZN(n27) );
  INV_X1 U64 ( .A(data_in[7]), .ZN(n65) );
  OAI22_X1 U65 ( .A1(n39), .A2(n64), .B1(net108202), .B2(n36), .ZN(n26) );
  INV_X1 U66 ( .A(data_in[8]), .ZN(n64) );
  OAI22_X1 U67 ( .A1(n40), .A2(n63), .B1(net108203), .B2(n36), .ZN(n25) );
  INV_X1 U68 ( .A(data_in[9]), .ZN(n63) );
  OAI22_X1 U69 ( .A1(n40), .A2(n62), .B1(net108204), .B2(n36), .ZN(n24) );
  INV_X1 U70 ( .A(data_in[10]), .ZN(n62) );
  OAI22_X1 U71 ( .A1(n40), .A2(n61), .B1(net108205), .B2(n36), .ZN(n23) );
  INV_X1 U72 ( .A(data_in[11]), .ZN(n61) );
  OAI22_X1 U73 ( .A1(n40), .A2(n60), .B1(net108206), .B2(n36), .ZN(n22) );
  INV_X1 U74 ( .A(data_in[12]), .ZN(n60) );
  NAND2_X1 U75 ( .A1(load), .A2(enable), .ZN(n90) );
  INV_X1 U76 ( .A(reset), .ZN(n3) );
  INV_X1 U77 ( .A(data_in[17]), .ZN(n54) );
  OAI22_X1 U78 ( .A1(n40), .A2(n59), .B1(net108207), .B2(n36), .ZN(n21) );
  INV_X1 U79 ( .A(data_in[20]), .ZN(n51) );
  INV_X1 U80 ( .A(data_in[16]), .ZN(n55) );
endmodule


module NRegister_N32_113 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, net108194, net108195, net108196, net108197,
         net108198, net108199, net108200, net108201, net108202, net108203,
         net108204, net108205, net108206, net108207, net108208, net108209,
         net108210, net108211, net108212, net108213, net108214, net108215,
         net108216, net108217, net108218, net108219, net108220, net108221,
         net108222, net108223, net108224, net108225, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n70, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n44), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n44), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n44), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n46), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n44), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n46), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n46), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n46), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n44), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n46), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n46), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n46), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n46), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n45), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n45), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n45), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n45), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n45), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n45), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n45), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n45), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n45), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n44), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n44), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n44), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n44), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n44), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n44), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n44), .Q(data_out[0]), 
        .QN(net108194) );
  INV_X1 U3 ( .A(n43), .ZN(n36) );
  INV_X1 U4 ( .A(n43), .ZN(n35) );
  BUF_X1 U5 ( .A(n90), .Z(n39) );
  BUF_X1 U6 ( .A(n90), .Z(n40) );
  BUF_X1 U7 ( .A(n90), .Z(n42) );
  BUF_X1 U8 ( .A(n90), .Z(n37) );
  BUF_X1 U9 ( .A(n90), .Z(n38) );
  BUF_X1 U10 ( .A(n90), .Z(n41) );
  BUF_X1 U11 ( .A(n90), .Z(n43) );
  BUF_X1 U12 ( .A(n3), .Z(n45) );
  BUF_X1 U13 ( .A(n3), .Z(n44) );
  BUF_X1 U14 ( .A(n3), .Z(n46) );
  OAI22_X1 U15 ( .A1(n38), .A2(n83), .B1(net108194), .B2(n36), .ZN(n34) );
  INV_X1 U16 ( .A(data_in[0]), .ZN(n83) );
  OAI22_X1 U17 ( .A1(n38), .A2(n82), .B1(net108195), .B2(n35), .ZN(n33) );
  INV_X1 U18 ( .A(data_in[1]), .ZN(n82) );
  OAI22_X1 U19 ( .A1(n37), .A2(n89), .B1(net108219), .B2(n36), .ZN(n9) );
  INV_X1 U20 ( .A(data_in[25]), .ZN(n89) );
  OAI22_X1 U21 ( .A1(n37), .A2(n88), .B1(net108220), .B2(n35), .ZN(n8) );
  INV_X1 U22 ( .A(data_in[26]), .ZN(n88) );
  OAI22_X1 U23 ( .A1(n37), .A2(n87), .B1(net108221), .B2(n36), .ZN(n7) );
  INV_X1 U24 ( .A(data_in[27]), .ZN(n87) );
  OAI22_X1 U25 ( .A1(n37), .A2(n86), .B1(net108222), .B2(n35), .ZN(n6) );
  INV_X1 U26 ( .A(data_in[28]), .ZN(n86) );
  OAI22_X1 U27 ( .A1(n37), .A2(n85), .B1(net108223), .B2(n36), .ZN(n5) );
  INV_X1 U28 ( .A(data_in[29]), .ZN(n85) );
  OAI22_X1 U29 ( .A1(n38), .A2(n84), .B1(net108224), .B2(n35), .ZN(n4) );
  INV_X1 U30 ( .A(data_in[30]), .ZN(n84) );
  OAI22_X1 U31 ( .A1(n38), .A2(n81), .B1(net108196), .B2(n36), .ZN(n32) );
  INV_X1 U32 ( .A(data_in[2]), .ZN(n81) );
  OAI22_X1 U33 ( .A1(n38), .A2(n80), .B1(net108197), .B2(n36), .ZN(n31) );
  INV_X1 U34 ( .A(data_in[3]), .ZN(n80) );
  OAI22_X1 U35 ( .A1(n39), .A2(n70), .B1(net108198), .B2(n36), .ZN(n30) );
  INV_X1 U36 ( .A(data_in[4]), .ZN(n70) );
  OAI22_X1 U37 ( .A1(n39), .A2(n67), .B1(net108199), .B2(n36), .ZN(n29) );
  INV_X1 U38 ( .A(data_in[5]), .ZN(n67) );
  OAI22_X1 U39 ( .A1(n39), .A2(n66), .B1(net108200), .B2(n36), .ZN(n28) );
  INV_X1 U40 ( .A(data_in[6]), .ZN(n66) );
  OAI22_X1 U41 ( .A1(n39), .A2(n65), .B1(net108201), .B2(n36), .ZN(n27) );
  INV_X1 U42 ( .A(data_in[7]), .ZN(n65) );
  OAI22_X1 U43 ( .A1(n39), .A2(n64), .B1(net108202), .B2(n36), .ZN(n26) );
  INV_X1 U44 ( .A(data_in[8]), .ZN(n64) );
  OAI22_X1 U45 ( .A1(n40), .A2(n63), .B1(net108203), .B2(n36), .ZN(n25) );
  INV_X1 U46 ( .A(data_in[9]), .ZN(n63) );
  OAI22_X1 U47 ( .A1(n40), .A2(n62), .B1(net108204), .B2(n36), .ZN(n24) );
  INV_X1 U48 ( .A(data_in[10]), .ZN(n62) );
  OAI22_X1 U49 ( .A1(n40), .A2(n61), .B1(net108205), .B2(n36), .ZN(n23) );
  INV_X1 U50 ( .A(data_in[11]), .ZN(n61) );
  OAI22_X1 U51 ( .A1(n40), .A2(n60), .B1(net108206), .B2(n36), .ZN(n22) );
  INV_X1 U52 ( .A(data_in[12]), .ZN(n60) );
  OAI22_X1 U53 ( .A1(n40), .A2(n59), .B1(net108207), .B2(n36), .ZN(n21) );
  INV_X1 U54 ( .A(data_in[13]), .ZN(n59) );
  OAI22_X1 U55 ( .A1(n41), .A2(n58), .B1(net108208), .B2(n35), .ZN(n20) );
  INV_X1 U56 ( .A(data_in[14]), .ZN(n58) );
  OAI22_X1 U57 ( .A1(n41), .A2(n56), .B1(net108209), .B2(n35), .ZN(n19) );
  INV_X1 U58 ( .A(data_in[15]), .ZN(n56) );
  OAI22_X1 U59 ( .A1(n41), .A2(n55), .B1(net108210), .B2(n35), .ZN(n18) );
  INV_X1 U60 ( .A(data_in[16]), .ZN(n55) );
  OAI22_X1 U61 ( .A1(n41), .A2(n54), .B1(net108211), .B2(n35), .ZN(n17) );
  INV_X1 U62 ( .A(data_in[17]), .ZN(n54) );
  OAI22_X1 U63 ( .A1(n42), .A2(n53), .B1(net108212), .B2(n35), .ZN(n16) );
  INV_X1 U64 ( .A(data_in[18]), .ZN(n53) );
  OAI22_X1 U65 ( .A1(n42), .A2(n52), .B1(net108213), .B2(n35), .ZN(n15) );
  INV_X1 U66 ( .A(data_in[19]), .ZN(n52) );
  OAI22_X1 U67 ( .A1(n42), .A2(n51), .B1(net108214), .B2(n35), .ZN(n14) );
  INV_X1 U68 ( .A(data_in[20]), .ZN(n51) );
  OAI22_X1 U69 ( .A1(n42), .A2(n50), .B1(net108215), .B2(n35), .ZN(n13) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n50) );
  OAI22_X1 U71 ( .A1(n42), .A2(n49), .B1(net108216), .B2(n35), .ZN(n12) );
  INV_X1 U72 ( .A(data_in[22]), .ZN(n49) );
  OAI22_X1 U73 ( .A1(n43), .A2(n48), .B1(net108217), .B2(n35), .ZN(n11) );
  INV_X1 U74 ( .A(data_in[23]), .ZN(n48) );
  OAI22_X1 U75 ( .A1(n43), .A2(n47), .B1(net108218), .B2(n35), .ZN(n10) );
  INV_X1 U76 ( .A(data_in[24]), .ZN(n47) );
  OAI22_X1 U77 ( .A1(n41), .A2(n57), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U78 ( .A(data_in[31]), .ZN(n57) );
  NAND2_X1 U79 ( .A1(load), .A2(enable), .ZN(n90) );
  INV_X1 U80 ( .A(reset), .ZN(n3) );
endmodule


module NRegister_N32_112 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, net108194, net108195, net108196, net108197,
         net108198, net108199, net108200, net108201, net108202, net108203,
         net108204, net108205, net108206, net108207, net108208, net108209,
         net108210, net108211, net108212, net108213, net108214, net108215,
         net108216, net108217, net108218, net108219, net108220, net108221,
         net108222, net108223, net108224, net108225, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n70, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n44), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n44), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n44), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n46), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n44), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n46), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n46), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n46), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n44), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n46), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n46), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n46), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n46), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n45), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n45), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n45), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n45), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n45), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n45), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n45), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n45), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n45), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n44), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n44), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n44), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n44), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n44), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n44), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n44), .Q(data_out[0]), 
        .QN(net108194) );
  INV_X1 U3 ( .A(n43), .ZN(n36) );
  INV_X1 U4 ( .A(n43), .ZN(n35) );
  BUF_X1 U5 ( .A(n90), .Z(n39) );
  BUF_X1 U6 ( .A(n90), .Z(n40) );
  BUF_X1 U7 ( .A(n90), .Z(n42) );
  BUF_X1 U8 ( .A(n90), .Z(n37) );
  BUF_X1 U9 ( .A(n90), .Z(n38) );
  BUF_X1 U10 ( .A(n90), .Z(n41) );
  BUF_X1 U11 ( .A(n90), .Z(n43) );
  BUF_X1 U12 ( .A(n3), .Z(n45) );
  BUF_X1 U13 ( .A(n3), .Z(n44) );
  BUF_X1 U14 ( .A(n3), .Z(n46) );
  OAI22_X1 U15 ( .A1(n38), .A2(n83), .B1(net108194), .B2(n36), .ZN(n34) );
  INV_X1 U16 ( .A(data_in[0]), .ZN(n83) );
  OAI22_X1 U17 ( .A1(n37), .A2(n86), .B1(net108222), .B2(n35), .ZN(n6) );
  INV_X1 U18 ( .A(data_in[28]), .ZN(n86) );
  OAI22_X1 U19 ( .A1(n38), .A2(n84), .B1(net108224), .B2(n36), .ZN(n4) );
  INV_X1 U20 ( .A(data_in[30]), .ZN(n84) );
  OAI22_X1 U21 ( .A1(n39), .A2(n64), .B1(net108202), .B2(n36), .ZN(n26) );
  INV_X1 U22 ( .A(data_in[8]), .ZN(n64) );
  OAI22_X1 U23 ( .A1(n40), .A2(n61), .B1(net108205), .B2(n36), .ZN(n23) );
  INV_X1 U24 ( .A(data_in[11]), .ZN(n61) );
  OAI22_X1 U25 ( .A1(n40), .A2(n59), .B1(net108207), .B2(n36), .ZN(n21) );
  INV_X1 U26 ( .A(data_in[13]), .ZN(n59) );
  OAI22_X1 U27 ( .A1(n41), .A2(n55), .B1(net108210), .B2(n35), .ZN(n18) );
  INV_X1 U28 ( .A(data_in[16]), .ZN(n55) );
  OAI22_X1 U29 ( .A1(n41), .A2(n54), .B1(net108211), .B2(n35), .ZN(n17) );
  INV_X1 U30 ( .A(data_in[17]), .ZN(n54) );
  OAI22_X1 U31 ( .A1(n42), .A2(n53), .B1(net108212), .B2(n35), .ZN(n16) );
  INV_X1 U32 ( .A(data_in[18]), .ZN(n53) );
  OAI22_X1 U33 ( .A1(n42), .A2(n52), .B1(net108213), .B2(n35), .ZN(n15) );
  INV_X1 U34 ( .A(data_in[19]), .ZN(n52) );
  OAI22_X1 U35 ( .A1(n42), .A2(n51), .B1(net108214), .B2(n35), .ZN(n14) );
  INV_X1 U36 ( .A(data_in[20]), .ZN(n51) );
  OAI22_X1 U37 ( .A1(n42), .A2(n49), .B1(net108216), .B2(n35), .ZN(n12) );
  INV_X1 U38 ( .A(data_in[22]), .ZN(n49) );
  OAI22_X1 U39 ( .A1(n43), .A2(n48), .B1(net108217), .B2(n35), .ZN(n11) );
  INV_X1 U40 ( .A(data_in[23]), .ZN(n48) );
  NAND2_X1 U41 ( .A1(load), .A2(enable), .ZN(n90) );
  OAI22_X1 U42 ( .A1(n38), .A2(n82), .B1(net108195), .B2(n35), .ZN(n33) );
  INV_X1 U43 ( .A(data_in[1]), .ZN(n82) );
  OAI22_X1 U44 ( .A1(n40), .A2(n63), .B1(net108203), .B2(n36), .ZN(n25) );
  INV_X1 U45 ( .A(data_in[9]), .ZN(n63) );
  OAI22_X1 U46 ( .A1(n40), .A2(n62), .B1(net108204), .B2(n36), .ZN(n24) );
  INV_X1 U47 ( .A(data_in[10]), .ZN(n62) );
  OAI22_X1 U48 ( .A1(n40), .A2(n60), .B1(net108206), .B2(n36), .ZN(n22) );
  INV_X1 U49 ( .A(data_in[12]), .ZN(n60) );
  OAI22_X1 U50 ( .A1(n41), .A2(n58), .B1(net108208), .B2(n35), .ZN(n20) );
  INV_X1 U51 ( .A(data_in[14]), .ZN(n58) );
  OAI22_X1 U52 ( .A1(n41), .A2(n56), .B1(net108209), .B2(n35), .ZN(n19) );
  INV_X1 U53 ( .A(data_in[15]), .ZN(n56) );
  OAI22_X1 U54 ( .A1(n42), .A2(n50), .B1(net108215), .B2(n35), .ZN(n13) );
  INV_X1 U55 ( .A(data_in[21]), .ZN(n50) );
  OAI22_X1 U56 ( .A1(n43), .A2(n47), .B1(net108218), .B2(n35), .ZN(n10) );
  INV_X1 U57 ( .A(data_in[24]), .ZN(n47) );
  OAI22_X1 U58 ( .A1(n37), .A2(n89), .B1(net108219), .B2(n36), .ZN(n9) );
  INV_X1 U59 ( .A(data_in[25]), .ZN(n89) );
  OAI22_X1 U60 ( .A1(n37), .A2(n88), .B1(net108220), .B2(n35), .ZN(n8) );
  INV_X1 U61 ( .A(data_in[26]), .ZN(n88) );
  OAI22_X1 U62 ( .A1(n37), .A2(n87), .B1(net108221), .B2(n36), .ZN(n7) );
  INV_X1 U63 ( .A(data_in[27]), .ZN(n87) );
  OAI22_X1 U64 ( .A1(n37), .A2(n85), .B1(net108223), .B2(n35), .ZN(n5) );
  INV_X1 U65 ( .A(data_in[29]), .ZN(n85) );
  OAI22_X1 U66 ( .A1(n39), .A2(n65), .B1(net108201), .B2(n36), .ZN(n27) );
  INV_X1 U67 ( .A(data_in[7]), .ZN(n65) );
  OAI22_X1 U68 ( .A1(n38), .A2(n81), .B1(net108196), .B2(n36), .ZN(n32) );
  INV_X1 U69 ( .A(data_in[2]), .ZN(n81) );
  OAI22_X1 U70 ( .A1(n38), .A2(n80), .B1(net108197), .B2(n36), .ZN(n31) );
  INV_X1 U71 ( .A(data_in[3]), .ZN(n80) );
  OAI22_X1 U72 ( .A1(n39), .A2(n70), .B1(net108198), .B2(n36), .ZN(n30) );
  INV_X1 U73 ( .A(data_in[4]), .ZN(n70) );
  OAI22_X1 U74 ( .A1(n39), .A2(n67), .B1(net108199), .B2(n36), .ZN(n29) );
  INV_X1 U75 ( .A(data_in[5]), .ZN(n67) );
  OAI22_X1 U76 ( .A1(n39), .A2(n66), .B1(net108200), .B2(n36), .ZN(n28) );
  INV_X1 U77 ( .A(data_in[6]), .ZN(n66) );
  OAI22_X1 U78 ( .A1(n41), .A2(n57), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U79 ( .A(data_in[31]), .ZN(n57) );
  INV_X1 U80 ( .A(reset), .ZN(n3) );
endmodule


module NRegister_N32_111 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, net108194, net108195, net108196, net108197,
         net108198, net108199, net108200, net108201, net108202, net108203,
         net108204, net108205, net108206, net108207, net108208, net108209,
         net108210, net108211, net108212, net108213, net108214, net108215,
         net108216, net108217, net108218, net108219, net108220, net108221,
         net108222, net108223, net108224, net108225, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n70, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n44), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n44), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n44), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n46), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n44), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n46), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n46), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n46), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n44), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n46), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n46), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n46), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n46), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n45), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n45), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n45), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n45), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n45), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n45), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n45), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n45), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n45), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n44), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n44), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n44), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n44), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n44), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n44), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n44), .Q(data_out[0]), 
        .QN(net108194) );
  INV_X1 U3 ( .A(n43), .ZN(n36) );
  INV_X1 U4 ( .A(n43), .ZN(n35) );
  BUF_X1 U5 ( .A(n90), .Z(n39) );
  BUF_X1 U6 ( .A(n90), .Z(n40) );
  BUF_X1 U7 ( .A(n90), .Z(n42) );
  BUF_X1 U8 ( .A(n90), .Z(n37) );
  BUF_X1 U9 ( .A(n90), .Z(n38) );
  BUF_X1 U10 ( .A(n90), .Z(n41) );
  BUF_X1 U11 ( .A(n90), .Z(n43) );
  BUF_X1 U12 ( .A(n3), .Z(n45) );
  BUF_X1 U13 ( .A(n3), .Z(n44) );
  BUF_X1 U14 ( .A(n3), .Z(n46) );
  OAI22_X1 U15 ( .A1(n38), .A2(n83), .B1(net108194), .B2(n36), .ZN(n34) );
  INV_X1 U16 ( .A(data_in[0]), .ZN(n83) );
  OAI22_X1 U17 ( .A1(n38), .A2(n82), .B1(net108195), .B2(n35), .ZN(n33) );
  INV_X1 U18 ( .A(data_in[1]), .ZN(n82) );
  OAI22_X1 U19 ( .A1(n37), .A2(n89), .B1(net108219), .B2(n36), .ZN(n9) );
  INV_X1 U20 ( .A(data_in[25]), .ZN(n89) );
  OAI22_X1 U21 ( .A1(n37), .A2(n88), .B1(net108220), .B2(n35), .ZN(n8) );
  INV_X1 U22 ( .A(data_in[26]), .ZN(n88) );
  OAI22_X1 U23 ( .A1(n37), .A2(n87), .B1(net108221), .B2(n36), .ZN(n7) );
  INV_X1 U24 ( .A(data_in[27]), .ZN(n87) );
  OAI22_X1 U25 ( .A1(n37), .A2(n86), .B1(net108222), .B2(n35), .ZN(n6) );
  INV_X1 U26 ( .A(data_in[28]), .ZN(n86) );
  OAI22_X1 U27 ( .A1(n37), .A2(n85), .B1(net108223), .B2(n36), .ZN(n5) );
  INV_X1 U28 ( .A(data_in[29]), .ZN(n85) );
  OAI22_X1 U29 ( .A1(n38), .A2(n84), .B1(net108224), .B2(n35), .ZN(n4) );
  INV_X1 U30 ( .A(data_in[30]), .ZN(n84) );
  OAI22_X1 U31 ( .A1(n38), .A2(n81), .B1(net108196), .B2(n36), .ZN(n32) );
  INV_X1 U32 ( .A(data_in[2]), .ZN(n81) );
  OAI22_X1 U33 ( .A1(n38), .A2(n80), .B1(net108197), .B2(n36), .ZN(n31) );
  INV_X1 U34 ( .A(data_in[3]), .ZN(n80) );
  OAI22_X1 U35 ( .A1(n39), .A2(n70), .B1(net108198), .B2(n36), .ZN(n30) );
  INV_X1 U36 ( .A(data_in[4]), .ZN(n70) );
  OAI22_X1 U37 ( .A1(n39), .A2(n67), .B1(net108199), .B2(n36), .ZN(n29) );
  INV_X1 U38 ( .A(data_in[5]), .ZN(n67) );
  OAI22_X1 U39 ( .A1(n39), .A2(n66), .B1(net108200), .B2(n36), .ZN(n28) );
  INV_X1 U40 ( .A(data_in[6]), .ZN(n66) );
  OAI22_X1 U41 ( .A1(n39), .A2(n65), .B1(net108201), .B2(n36), .ZN(n27) );
  INV_X1 U42 ( .A(data_in[7]), .ZN(n65) );
  OAI22_X1 U43 ( .A1(n39), .A2(n64), .B1(net108202), .B2(n36), .ZN(n26) );
  INV_X1 U44 ( .A(data_in[8]), .ZN(n64) );
  OAI22_X1 U45 ( .A1(n40), .A2(n63), .B1(net108203), .B2(n36), .ZN(n25) );
  INV_X1 U46 ( .A(data_in[9]), .ZN(n63) );
  OAI22_X1 U47 ( .A1(n40), .A2(n62), .B1(net108204), .B2(n36), .ZN(n24) );
  INV_X1 U48 ( .A(data_in[10]), .ZN(n62) );
  OAI22_X1 U49 ( .A1(n40), .A2(n61), .B1(net108205), .B2(n36), .ZN(n23) );
  OAI22_X1 U50 ( .A1(n40), .A2(n60), .B1(net108206), .B2(n36), .ZN(n22) );
  OAI22_X1 U51 ( .A1(n40), .A2(n59), .B1(net108207), .B2(n36), .ZN(n21) );
  OAI22_X1 U52 ( .A1(n41), .A2(n58), .B1(net108208), .B2(n35), .ZN(n20) );
  INV_X1 U53 ( .A(data_in[14]), .ZN(n58) );
  OAI22_X1 U54 ( .A1(n41), .A2(n56), .B1(net108209), .B2(n35), .ZN(n19) );
  OAI22_X1 U55 ( .A1(n41), .A2(n55), .B1(net108210), .B2(n35), .ZN(n18) );
  OAI22_X1 U56 ( .A1(n41), .A2(n54), .B1(net108211), .B2(n35), .ZN(n17) );
  OAI22_X1 U57 ( .A1(n42), .A2(n53), .B1(net108212), .B2(n35), .ZN(n16) );
  OAI22_X1 U58 ( .A1(n42), .A2(n52), .B1(net108213), .B2(n35), .ZN(n15) );
  OAI22_X1 U59 ( .A1(n42), .A2(n51), .B1(net108214), .B2(n35), .ZN(n14) );
  OAI22_X1 U60 ( .A1(n42), .A2(n50), .B1(net108215), .B2(n35), .ZN(n13) );
  INV_X1 U61 ( .A(data_in[21]), .ZN(n50) );
  OAI22_X1 U62 ( .A1(n42), .A2(n49), .B1(net108216), .B2(n35), .ZN(n12) );
  INV_X1 U63 ( .A(data_in[22]), .ZN(n49) );
  OAI22_X1 U64 ( .A1(n43), .A2(n48), .B1(net108217), .B2(n35), .ZN(n11) );
  INV_X1 U65 ( .A(data_in[23]), .ZN(n48) );
  OAI22_X1 U66 ( .A1(n43), .A2(n47), .B1(net108218), .B2(n35), .ZN(n10) );
  INV_X1 U67 ( .A(data_in[24]), .ZN(n47) );
  OAI22_X1 U68 ( .A1(n41), .A2(n57), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U69 ( .A(data_in[31]), .ZN(n57) );
  NAND2_X1 U70 ( .A1(load), .A2(enable), .ZN(n90) );
  INV_X1 U71 ( .A(reset), .ZN(n3) );
  INV_X1 U72 ( .A(data_in[13]), .ZN(n59) );
  INV_X1 U73 ( .A(data_in[15]), .ZN(n56) );
  INV_X1 U74 ( .A(data_in[16]), .ZN(n55) );
  INV_X1 U75 ( .A(data_in[18]), .ZN(n53) );
  INV_X1 U76 ( .A(data_in[17]), .ZN(n54) );
  INV_X1 U77 ( .A(data_in[19]), .ZN(n52) );
  INV_X1 U78 ( .A(data_in[11]), .ZN(n61) );
  INV_X1 U79 ( .A(data_in[20]), .ZN(n51) );
  INV_X1 U80 ( .A(data_in[12]), .ZN(n60) );
endmodule


module NRegister_N32_110 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108194, net108195, net108196, net108197, net108198,
         net108199, net108200, net108201, net108202, net108203, net108204,
         net108205, net108206, net108207, net108208, net108209, net108210,
         net108211, net108212, net108213, net108214, net108215, net108216,
         net108217, net108218, net108219, net108220, net108221, net108222,
         net108223, net108224, net108225, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n46), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n46), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n46), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n44), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n46), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n44), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n44), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n44), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n46), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n44), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n44), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n44), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n44), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n44), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n44), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n44), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n44), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n45), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n45), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n45), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n45), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n45), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n45), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n45), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n45), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n45), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n46), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n46), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n46), .Q(data_out[0]), 
        .QN(net108194) );
  INV_X1 U3 ( .A(n43), .ZN(n36) );
  INV_X1 U4 ( .A(n43), .ZN(n35) );
  BUF_X1 U5 ( .A(n92), .Z(n39) );
  BUF_X1 U6 ( .A(n92), .Z(n40) );
  BUF_X1 U7 ( .A(n92), .Z(n42) );
  BUF_X1 U8 ( .A(n92), .Z(n37) );
  BUF_X1 U9 ( .A(n92), .Z(n38) );
  BUF_X1 U10 ( .A(n92), .Z(n41) );
  BUF_X1 U11 ( .A(n92), .Z(n43) );
  BUF_X1 U12 ( .A(n47), .Z(n45) );
  BUF_X1 U13 ( .A(n47), .Z(n44) );
  BUF_X1 U14 ( .A(n47), .Z(n46) );
  OAI22_X1 U15 ( .A1(n38), .A2(n85), .B1(net108194), .B2(n36), .ZN(n34) );
  INV_X1 U16 ( .A(data_in[0]), .ZN(n85) );
  OAI22_X1 U17 ( .A1(n38), .A2(n84), .B1(net108195), .B2(n35), .ZN(n33) );
  INV_X1 U18 ( .A(data_in[1]), .ZN(n84) );
  OAI22_X1 U19 ( .A1(n37), .A2(n91), .B1(net108219), .B2(n36), .ZN(n9) );
  INV_X1 U20 ( .A(data_in[25]), .ZN(n91) );
  OAI22_X1 U21 ( .A1(n37), .A2(n90), .B1(net108220), .B2(n35), .ZN(n8) );
  INV_X1 U22 ( .A(data_in[26]), .ZN(n90) );
  OAI22_X1 U23 ( .A1(n37), .A2(n89), .B1(net108221), .B2(n36), .ZN(n7) );
  INV_X1 U24 ( .A(data_in[27]), .ZN(n89) );
  OAI22_X1 U25 ( .A1(n37), .A2(n88), .B1(net108222), .B2(n35), .ZN(n6) );
  INV_X1 U26 ( .A(data_in[28]), .ZN(n88) );
  OAI22_X1 U27 ( .A1(n37), .A2(n87), .B1(net108223), .B2(n36), .ZN(n5) );
  INV_X1 U28 ( .A(data_in[29]), .ZN(n87) );
  OAI22_X1 U29 ( .A1(n38), .A2(n86), .B1(net108224), .B2(n35), .ZN(n4) );
  INV_X1 U30 ( .A(data_in[30]), .ZN(n86) );
  OAI22_X1 U31 ( .A1(n38), .A2(n83), .B1(net108196), .B2(n36), .ZN(n32) );
  INV_X1 U32 ( .A(data_in[2]), .ZN(n83) );
  OAI22_X1 U33 ( .A1(n38), .A2(n82), .B1(net108197), .B2(n36), .ZN(n31) );
  INV_X1 U34 ( .A(data_in[3]), .ZN(n82) );
  OAI22_X1 U35 ( .A1(n39), .A2(n81), .B1(net108198), .B2(n36), .ZN(n30) );
  INV_X1 U36 ( .A(data_in[4]), .ZN(n81) );
  OAI22_X1 U37 ( .A1(n39), .A2(n70), .B1(net108199), .B2(n36), .ZN(n29) );
  INV_X1 U38 ( .A(data_in[5]), .ZN(n70) );
  OAI22_X1 U39 ( .A1(n39), .A2(n67), .B1(net108200), .B2(n36), .ZN(n28) );
  INV_X1 U40 ( .A(data_in[6]), .ZN(n67) );
  OAI22_X1 U41 ( .A1(n39), .A2(n66), .B1(net108201), .B2(n36), .ZN(n27) );
  INV_X1 U42 ( .A(data_in[7]), .ZN(n66) );
  OAI22_X1 U43 ( .A1(n39), .A2(n65), .B1(net108202), .B2(n36), .ZN(n26) );
  INV_X1 U44 ( .A(data_in[8]), .ZN(n65) );
  OAI22_X1 U45 ( .A1(n40), .A2(n64), .B1(net108203), .B2(n36), .ZN(n25) );
  INV_X1 U46 ( .A(data_in[9]), .ZN(n64) );
  OAI22_X1 U47 ( .A1(n40), .A2(n63), .B1(net108204), .B2(n36), .ZN(n24) );
  INV_X1 U48 ( .A(data_in[10]), .ZN(n63) );
  OAI22_X1 U49 ( .A1(n40), .A2(n62), .B1(net108205), .B2(n36), .ZN(n23) );
  INV_X1 U50 ( .A(data_in[11]), .ZN(n62) );
  OAI22_X1 U51 ( .A1(n40), .A2(n61), .B1(net108206), .B2(n36), .ZN(n22) );
  INV_X1 U52 ( .A(data_in[12]), .ZN(n61) );
  OAI22_X1 U53 ( .A1(n40), .A2(n60), .B1(net108207), .B2(n36), .ZN(n21) );
  INV_X1 U54 ( .A(data_in[13]), .ZN(n60) );
  OAI22_X1 U55 ( .A1(n41), .A2(n59), .B1(net108208), .B2(n35), .ZN(n20) );
  INV_X1 U56 ( .A(data_in[14]), .ZN(n59) );
  OAI22_X1 U57 ( .A1(n41), .A2(n57), .B1(net108209), .B2(n35), .ZN(n19) );
  INV_X1 U58 ( .A(data_in[15]), .ZN(n57) );
  OAI22_X1 U59 ( .A1(n41), .A2(n56), .B1(net108210), .B2(n35), .ZN(n18) );
  INV_X1 U60 ( .A(data_in[16]), .ZN(n56) );
  OAI22_X1 U61 ( .A1(n41), .A2(n55), .B1(net108211), .B2(n35), .ZN(n17) );
  INV_X1 U62 ( .A(data_in[17]), .ZN(n55) );
  OAI22_X1 U63 ( .A1(n42), .A2(n54), .B1(net108212), .B2(n35), .ZN(n16) );
  INV_X1 U64 ( .A(data_in[18]), .ZN(n54) );
  OAI22_X1 U65 ( .A1(n42), .A2(n53), .B1(net108213), .B2(n35), .ZN(n15) );
  INV_X1 U66 ( .A(data_in[19]), .ZN(n53) );
  OAI22_X1 U67 ( .A1(n42), .A2(n52), .B1(net108214), .B2(n35), .ZN(n14) );
  INV_X1 U68 ( .A(data_in[20]), .ZN(n52) );
  OAI22_X1 U69 ( .A1(n42), .A2(n51), .B1(net108215), .B2(n35), .ZN(n13) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n51) );
  OAI22_X1 U71 ( .A1(n42), .A2(n50), .B1(net108216), .B2(n35), .ZN(n12) );
  INV_X1 U72 ( .A(data_in[22]), .ZN(n50) );
  OAI22_X1 U73 ( .A1(n43), .A2(n49), .B1(net108217), .B2(n35), .ZN(n11) );
  INV_X1 U74 ( .A(data_in[23]), .ZN(n49) );
  OAI22_X1 U75 ( .A1(n43), .A2(n48), .B1(net108218), .B2(n35), .ZN(n10) );
  INV_X1 U76 ( .A(data_in[24]), .ZN(n48) );
  OAI22_X1 U77 ( .A1(n41), .A2(n58), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U78 ( .A(data_in[31]), .ZN(n58) );
  NAND2_X1 U79 ( .A1(load), .A2(enable), .ZN(n92) );
  INV_X1 U80 ( .A(reset), .ZN(n47) );
endmodule


module NRegister_N32_43 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108194, net108195, net108196, net108197, net108198,
         net108199, net108200, net108201, net108202, net108203, net108204,
         net108205, net108206, net108207, net108208, net108209, net108210,
         net108211, net108212, net108213, net108214, net108215, net108216,
         net108217, net108218, net108219, net108220, net108221, net108222,
         net108223, net108224, net108225, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n46), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n46), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n46), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n44), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n46), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n44), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n44), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n44), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n46), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n44), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n44), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n44), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n44), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n44), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n44), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n44), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n44), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n45), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n45), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n45), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n45), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n45), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n45), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n45), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n45), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n45), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n46), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n46), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n46), .Q(data_out[0]), 
        .QN(net108194) );
  BUF_X1 U3 ( .A(n47), .Z(n45) );
  BUF_X1 U4 ( .A(n47), .Z(n44) );
  BUF_X1 U5 ( .A(n47), .Z(n46) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n47) );
  BUF_X1 U9 ( .A(n92), .Z(n39) );
  BUF_X1 U10 ( .A(n92), .Z(n40) );
  BUF_X1 U11 ( .A(n92), .Z(n42) );
  BUF_X1 U12 ( .A(n92), .Z(n37) );
  BUF_X1 U13 ( .A(n92), .Z(n38) );
  BUF_X1 U14 ( .A(n92), .Z(n41) );
  BUF_X1 U15 ( .A(n92), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n84), .B1(net108195), .B2(n36), .ZN(n33) );
  INV_X1 U17 ( .A(data_in[1]), .ZN(n84) );
  OAI22_X1 U18 ( .A1(n37), .A2(n90), .B1(net108220), .B2(n35), .ZN(n8) );
  INV_X1 U19 ( .A(data_in[26]), .ZN(n90) );
  OAI22_X1 U20 ( .A1(n37), .A2(n89), .B1(net108221), .B2(n36), .ZN(n7) );
  INV_X1 U21 ( .A(data_in[27]), .ZN(n89) );
  OAI22_X1 U22 ( .A1(n37), .A2(n87), .B1(net108223), .B2(n35), .ZN(n5) );
  INV_X1 U23 ( .A(data_in[29]), .ZN(n87) );
  OAI22_X1 U24 ( .A1(n38), .A2(n83), .B1(net108196), .B2(n36), .ZN(n32) );
  INV_X1 U25 ( .A(data_in[2]), .ZN(n83) );
  OAI22_X1 U26 ( .A1(n38), .A2(n82), .B1(net108197), .B2(n36), .ZN(n31) );
  INV_X1 U27 ( .A(data_in[3]), .ZN(n82) );
  OAI22_X1 U28 ( .A1(n39), .A2(n81), .B1(net108198), .B2(n36), .ZN(n30) );
  INV_X1 U29 ( .A(data_in[4]), .ZN(n81) );
  OAI22_X1 U30 ( .A1(n39), .A2(n70), .B1(net108199), .B2(n36), .ZN(n29) );
  INV_X1 U31 ( .A(data_in[5]), .ZN(n70) );
  OAI22_X1 U32 ( .A1(n39), .A2(n67), .B1(net108200), .B2(n36), .ZN(n28) );
  INV_X1 U33 ( .A(data_in[6]), .ZN(n67) );
  OAI22_X1 U34 ( .A1(n40), .A2(n63), .B1(net108204), .B2(n36), .ZN(n24) );
  INV_X1 U35 ( .A(data_in[10]), .ZN(n63) );
  OAI22_X1 U36 ( .A1(n40), .A2(n62), .B1(net108205), .B2(n36), .ZN(n23) );
  INV_X1 U37 ( .A(data_in[11]), .ZN(n62) );
  OAI22_X1 U38 ( .A1(n41), .A2(n59), .B1(net108208), .B2(n35), .ZN(n20) );
  INV_X1 U39 ( .A(data_in[14]), .ZN(n59) );
  OAI22_X1 U40 ( .A1(n41), .A2(n57), .B1(net108209), .B2(n35), .ZN(n19) );
  INV_X1 U41 ( .A(data_in[15]), .ZN(n57) );
  OAI22_X1 U42 ( .A1(n41), .A2(n56), .B1(net108210), .B2(n35), .ZN(n18) );
  INV_X1 U43 ( .A(data_in[16]), .ZN(n56) );
  OAI22_X1 U44 ( .A1(n41), .A2(n55), .B1(net108211), .B2(n35), .ZN(n17) );
  INV_X1 U45 ( .A(data_in[17]), .ZN(n55) );
  OAI22_X1 U46 ( .A1(n42), .A2(n53), .B1(net108213), .B2(n35), .ZN(n15) );
  INV_X1 U47 ( .A(data_in[19]), .ZN(n53) );
  OAI22_X1 U48 ( .A1(n43), .A2(n49), .B1(net108217), .B2(n35), .ZN(n11) );
  INV_X1 U49 ( .A(data_in[23]), .ZN(n49) );
  OAI22_X1 U50 ( .A1(n43), .A2(n48), .B1(net108218), .B2(n35), .ZN(n10) );
  INV_X1 U51 ( .A(data_in[24]), .ZN(n48) );
  OAI22_X1 U52 ( .A1(n41), .A2(n58), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U53 ( .A(data_in[31]), .ZN(n58) );
  NAND2_X1 U54 ( .A1(load), .A2(enable), .ZN(n92) );
  OAI22_X1 U55 ( .A1(n38), .A2(n86), .B1(net108224), .B2(n36), .ZN(n4) );
  INV_X1 U56 ( .A(data_in[30]), .ZN(n86) );
  OAI22_X1 U57 ( .A1(n40), .A2(n64), .B1(net108203), .B2(n36), .ZN(n25) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n64) );
  OAI22_X1 U59 ( .A1(n39), .A2(n65), .B1(net108202), .B2(n36), .ZN(n26) );
  INV_X1 U60 ( .A(data_in[8]), .ZN(n65) );
  OAI22_X1 U61 ( .A1(n37), .A2(n91), .B1(net108219), .B2(n35), .ZN(n9) );
  INV_X1 U62 ( .A(data_in[25]), .ZN(n91) );
  OAI22_X1 U63 ( .A1(n42), .A2(n50), .B1(net108216), .B2(n35), .ZN(n12) );
  INV_X1 U64 ( .A(data_in[22]), .ZN(n50) );
  OAI22_X1 U65 ( .A1(n42), .A2(n51), .B1(net108215), .B2(n35), .ZN(n13) );
  INV_X1 U66 ( .A(data_in[21]), .ZN(n51) );
  OAI22_X1 U67 ( .A1(n42), .A2(n52), .B1(net108214), .B2(n35), .ZN(n14) );
  INV_X1 U68 ( .A(data_in[20]), .ZN(n52) );
  OAI22_X1 U69 ( .A1(n39), .A2(n66), .B1(net108201), .B2(n36), .ZN(n27) );
  INV_X1 U70 ( .A(data_in[7]), .ZN(n66) );
  OAI22_X1 U71 ( .A1(n37), .A2(n88), .B1(net108222), .B2(n36), .ZN(n6) );
  INV_X1 U72 ( .A(data_in[28]), .ZN(n88) );
  OAI22_X1 U73 ( .A1(n42), .A2(n54), .B1(net108212), .B2(n35), .ZN(n16) );
  INV_X1 U74 ( .A(data_in[18]), .ZN(n54) );
  OAI22_X1 U75 ( .A1(n40), .A2(n60), .B1(net108207), .B2(n36), .ZN(n21) );
  INV_X1 U76 ( .A(data_in[13]), .ZN(n60) );
  OAI22_X1 U77 ( .A1(n40), .A2(n61), .B1(net108206), .B2(n36), .ZN(n22) );
  INV_X1 U78 ( .A(data_in[12]), .ZN(n61) );
  OAI22_X1 U79 ( .A1(n38), .A2(n85), .B1(net108194), .B2(n35), .ZN(n34) );
  INV_X1 U80 ( .A(data_in[0]), .ZN(n85) );
endmodule


module NRegister_N32_42 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, net108194, net108195, net108196, net108197,
         net108198, net108199, net108200, net108201, net108202, net108203,
         net108204, net108205, net108206, net108207, net108208, net108209,
         net108210, net108211, net108212, net108213, net108214, net108215,
         net108216, net108217, net108218, net108219, net108220, net108221,
         net108222, net108223, net108224, net108225, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n70, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n44), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n44), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n44), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n46), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n44), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n46), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n46), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n46), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n44), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n46), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n46), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n46), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n46), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n45), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n45), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n45), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n45), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n45), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n45), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n45), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n45), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n45), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n44), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n44), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n44), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n44), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n44), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n44), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n44), .Q(data_out[0]), 
        .QN(net108194) );
  BUF_X1 U3 ( .A(n3), .Z(n45) );
  BUF_X1 U4 ( .A(n3), .Z(n44) );
  BUF_X1 U5 ( .A(n3), .Z(n46) );
  INV_X1 U6 ( .A(reset), .ZN(n3) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  BUF_X1 U8 ( .A(n90), .Z(n39) );
  BUF_X1 U9 ( .A(n90), .Z(n40) );
  BUF_X1 U10 ( .A(n90), .Z(n42) );
  BUF_X1 U11 ( .A(n90), .Z(n37) );
  BUF_X1 U12 ( .A(n90), .Z(n38) );
  BUF_X1 U13 ( .A(n90), .Z(n43) );
  BUF_X1 U14 ( .A(n90), .Z(n41) );
  OAI22_X1 U15 ( .A1(n37), .A2(n85), .B1(net108223), .B2(n36), .ZN(n5) );
  INV_X1 U16 ( .A(data_in[29]), .ZN(n85) );
  OAI22_X1 U17 ( .A1(n37), .A2(n86), .B1(net108222), .B2(n36), .ZN(n6) );
  INV_X1 U18 ( .A(data_in[28]), .ZN(n86) );
  OAI22_X1 U19 ( .A1(n37), .A2(n87), .B1(net108221), .B2(n36), .ZN(n7) );
  INV_X1 U20 ( .A(data_in[27]), .ZN(n87) );
  OAI22_X1 U21 ( .A1(n37), .A2(n88), .B1(net108220), .B2(n36), .ZN(n8) );
  INV_X1 U22 ( .A(data_in[26]), .ZN(n88) );
  OAI22_X1 U23 ( .A1(n38), .A2(n84), .B1(net108224), .B2(n36), .ZN(n4) );
  INV_X1 U24 ( .A(data_in[30]), .ZN(n84) );
  OAI22_X1 U25 ( .A1(n37), .A2(n89), .B1(net108219), .B2(n36), .ZN(n9) );
  INV_X1 U26 ( .A(data_in[25]), .ZN(n89) );
  OAI22_X1 U27 ( .A1(n38), .A2(n83), .B1(net108194), .B2(n36), .ZN(n34) );
  INV_X1 U28 ( .A(data_in[0]), .ZN(n83) );
  OAI22_X1 U29 ( .A1(n38), .A2(n82), .B1(net108195), .B2(n36), .ZN(n33) );
  INV_X1 U30 ( .A(data_in[1]), .ZN(n82) );
  OAI22_X1 U31 ( .A1(n40), .A2(n60), .B1(net108206), .B2(n35), .ZN(n22) );
  INV_X1 U32 ( .A(data_in[12]), .ZN(n60) );
  OAI22_X1 U33 ( .A1(n40), .A2(n59), .B1(net108207), .B2(n36), .ZN(n21) );
  INV_X1 U34 ( .A(data_in[13]), .ZN(n59) );
  OAI22_X1 U35 ( .A1(n39), .A2(n64), .B1(net108202), .B2(n35), .ZN(n26) );
  INV_X1 U36 ( .A(data_in[8]), .ZN(n64) );
  OAI22_X1 U37 ( .A1(n40), .A2(n63), .B1(net108203), .B2(n36), .ZN(n25) );
  INV_X1 U38 ( .A(data_in[9]), .ZN(n63) );
  OAI22_X1 U39 ( .A1(n40), .A2(n62), .B1(net108204), .B2(n35), .ZN(n24) );
  INV_X1 U40 ( .A(data_in[10]), .ZN(n62) );
  OAI22_X1 U41 ( .A1(n40), .A2(n61), .B1(net108205), .B2(n36), .ZN(n23) );
  INV_X1 U42 ( .A(data_in[11]), .ZN(n61) );
  OAI22_X1 U43 ( .A1(n43), .A2(n47), .B1(net108218), .B2(n35), .ZN(n10) );
  INV_X1 U44 ( .A(data_in[24]), .ZN(n47) );
  OAI22_X1 U45 ( .A1(n43), .A2(n48), .B1(net108217), .B2(n35), .ZN(n11) );
  INV_X1 U46 ( .A(data_in[23]), .ZN(n48) );
  OAI22_X1 U47 ( .A1(n42), .A2(n49), .B1(net108216), .B2(n35), .ZN(n12) );
  INV_X1 U48 ( .A(data_in[22]), .ZN(n49) );
  OAI22_X1 U49 ( .A1(n42), .A2(n50), .B1(net108215), .B2(n35), .ZN(n13) );
  INV_X1 U50 ( .A(data_in[21]), .ZN(n50) );
  OAI22_X1 U51 ( .A1(n42), .A2(n51), .B1(net108214), .B2(n35), .ZN(n14) );
  INV_X1 U52 ( .A(data_in[20]), .ZN(n51) );
  OAI22_X1 U53 ( .A1(n42), .A2(n52), .B1(net108213), .B2(n35), .ZN(n15) );
  INV_X1 U54 ( .A(data_in[19]), .ZN(n52) );
  OAI22_X1 U55 ( .A1(n42), .A2(n53), .B1(net108212), .B2(n35), .ZN(n16) );
  INV_X1 U56 ( .A(data_in[18]), .ZN(n53) );
  OAI22_X1 U57 ( .A1(n41), .A2(n58), .B1(net108208), .B2(n35), .ZN(n20) );
  INV_X1 U58 ( .A(data_in[14]), .ZN(n58) );
  OAI22_X1 U59 ( .A1(n41), .A2(n54), .B1(net108211), .B2(n35), .ZN(n17) );
  INV_X1 U60 ( .A(data_in[17]), .ZN(n54) );
  OAI22_X1 U61 ( .A1(n41), .A2(n55), .B1(net108210), .B2(n35), .ZN(n18) );
  INV_X1 U62 ( .A(data_in[16]), .ZN(n55) );
  OAI22_X1 U63 ( .A1(n41), .A2(n56), .B1(net108209), .B2(n35), .ZN(n19) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n56) );
  OAI22_X1 U65 ( .A1(n38), .A2(n81), .B1(net108196), .B2(n35), .ZN(n32) );
  INV_X1 U66 ( .A(data_in[2]), .ZN(n81) );
  OAI22_X1 U67 ( .A1(n38), .A2(n80), .B1(net108197), .B2(n36), .ZN(n31) );
  INV_X1 U68 ( .A(data_in[3]), .ZN(n80) );
  OAI22_X1 U69 ( .A1(n39), .A2(n70), .B1(net108198), .B2(n36), .ZN(n30) );
  INV_X1 U70 ( .A(data_in[4]), .ZN(n70) );
  OAI22_X1 U71 ( .A1(n39), .A2(n67), .B1(net108199), .B2(n36), .ZN(n29) );
  INV_X1 U72 ( .A(data_in[5]), .ZN(n67) );
  OAI22_X1 U73 ( .A1(n39), .A2(n66), .B1(net108200), .B2(n36), .ZN(n28) );
  INV_X1 U74 ( .A(data_in[6]), .ZN(n66) );
  OAI22_X1 U75 ( .A1(n39), .A2(n65), .B1(net108201), .B2(n36), .ZN(n27) );
  INV_X1 U76 ( .A(data_in[7]), .ZN(n65) );
  NAND2_X1 U77 ( .A1(load), .A2(enable), .ZN(n90) );
  OAI22_X1 U78 ( .A1(n57), .A2(n41), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U79 ( .A(data_in[31]), .ZN(n57) );
  INV_X1 U80 ( .A(n43), .ZN(n36) );
endmodule


module NRegister_N32_40 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, net108194, net108195, net108196, net108197,
         net108198, net108199, net108200, net108201, net108202, net108203,
         net108204, net108205, net108206, net108207, net108208, net108209,
         net108210, net108211, net108212, net108213, net108214, net108215,
         net108216, net108217, net108218, net108219, net108220, net108221,
         net108222, net108223, net108224, net108225, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n70, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n44), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n44), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n44), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n46), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n44), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n46), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n46), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n46), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n44), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n46), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n46), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n46), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n46), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n45), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n45), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n45), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n45), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n45), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n45), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n45), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n45), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n45), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n44), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n44), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n44), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n44), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n44), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n44), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n44), .Q(data_out[0]), 
        .QN(net108194) );
  BUF_X1 U3 ( .A(n3), .Z(n45) );
  BUF_X1 U4 ( .A(n3), .Z(n44) );
  BUF_X1 U5 ( .A(n3), .Z(n46) );
  INV_X1 U6 ( .A(reset), .ZN(n3) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n90), .Z(n39) );
  BUF_X1 U10 ( .A(n90), .Z(n40) );
  BUF_X1 U11 ( .A(n90), .Z(n42) );
  BUF_X1 U12 ( .A(n90), .Z(n37) );
  BUF_X1 U13 ( .A(n90), .Z(n38) );
  BUF_X1 U14 ( .A(n90), .Z(n41) );
  BUF_X1 U15 ( .A(n90), .Z(n43) );
  OAI22_X1 U16 ( .A1(n43), .A2(n48), .B1(net108217), .B2(n35), .ZN(n11) );
  INV_X1 U17 ( .A(data_in[23]), .ZN(n48) );
  OAI22_X1 U18 ( .A1(n43), .A2(n47), .B1(net108218), .B2(n35), .ZN(n10) );
  INV_X1 U19 ( .A(data_in[24]), .ZN(n47) );
  OAI22_X1 U20 ( .A1(n37), .A2(n89), .B1(net108219), .B2(n36), .ZN(n9) );
  INV_X1 U21 ( .A(data_in[25]), .ZN(n89) );
  OAI22_X1 U22 ( .A1(n37), .A2(n88), .B1(net108220), .B2(n35), .ZN(n8) );
  INV_X1 U23 ( .A(data_in[26]), .ZN(n88) );
  OAI22_X1 U24 ( .A1(n37), .A2(n87), .B1(net108221), .B2(n36), .ZN(n7) );
  INV_X1 U25 ( .A(data_in[27]), .ZN(n87) );
  OAI22_X1 U26 ( .A1(n37), .A2(n86), .B1(net108222), .B2(n35), .ZN(n6) );
  INV_X1 U27 ( .A(data_in[28]), .ZN(n86) );
  OAI22_X1 U28 ( .A1(n37), .A2(n85), .B1(net108223), .B2(n36), .ZN(n5) );
  INV_X1 U29 ( .A(data_in[29]), .ZN(n85) );
  OAI22_X1 U30 ( .A1(n38), .A2(n84), .B1(net108224), .B2(n35), .ZN(n4) );
  INV_X1 U31 ( .A(data_in[30]), .ZN(n84) );
  OAI22_X1 U32 ( .A1(n41), .A2(n57), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U33 ( .A(data_in[31]), .ZN(n57) );
  OAI22_X1 U34 ( .A1(n40), .A2(n60), .B1(net108206), .B2(n36), .ZN(n22) );
  INV_X1 U35 ( .A(data_in[12]), .ZN(n60) );
  OAI22_X1 U36 ( .A1(n40), .A2(n59), .B1(net108207), .B2(n36), .ZN(n21) );
  INV_X1 U37 ( .A(data_in[13]), .ZN(n59) );
  OAI22_X1 U38 ( .A1(n41), .A2(n58), .B1(net108208), .B2(n35), .ZN(n20) );
  INV_X1 U39 ( .A(data_in[14]), .ZN(n58) );
  OAI22_X1 U40 ( .A1(n41), .A2(n56), .B1(net108209), .B2(n35), .ZN(n19) );
  INV_X1 U41 ( .A(data_in[15]), .ZN(n56) );
  OAI22_X1 U42 ( .A1(n41), .A2(n55), .B1(net108210), .B2(n35), .ZN(n18) );
  INV_X1 U43 ( .A(data_in[16]), .ZN(n55) );
  OAI22_X1 U44 ( .A1(n41), .A2(n54), .B1(net108211), .B2(n35), .ZN(n17) );
  INV_X1 U45 ( .A(data_in[17]), .ZN(n54) );
  OAI22_X1 U46 ( .A1(n42), .A2(n53), .B1(net108212), .B2(n35), .ZN(n16) );
  INV_X1 U47 ( .A(data_in[18]), .ZN(n53) );
  OAI22_X1 U48 ( .A1(n42), .A2(n52), .B1(net108213), .B2(n35), .ZN(n15) );
  INV_X1 U49 ( .A(data_in[19]), .ZN(n52) );
  OAI22_X1 U50 ( .A1(n42), .A2(n51), .B1(net108214), .B2(n35), .ZN(n14) );
  INV_X1 U51 ( .A(data_in[20]), .ZN(n51) );
  OAI22_X1 U52 ( .A1(n42), .A2(n50), .B1(net108215), .B2(n35), .ZN(n13) );
  INV_X1 U53 ( .A(data_in[21]), .ZN(n50) );
  OAI22_X1 U54 ( .A1(n42), .A2(n49), .B1(net108216), .B2(n35), .ZN(n12) );
  INV_X1 U55 ( .A(data_in[22]), .ZN(n49) );
  OAI22_X1 U56 ( .A1(n38), .A2(n83), .B1(net108194), .B2(n36), .ZN(n34) );
  INV_X1 U57 ( .A(data_in[0]), .ZN(n83) );
  OAI22_X1 U58 ( .A1(n38), .A2(n82), .B1(net108195), .B2(n35), .ZN(n33) );
  INV_X1 U59 ( .A(data_in[1]), .ZN(n82) );
  OAI22_X1 U60 ( .A1(n38), .A2(n81), .B1(net108196), .B2(n36), .ZN(n32) );
  INV_X1 U61 ( .A(data_in[2]), .ZN(n81) );
  NAND2_X1 U62 ( .A1(load), .A2(enable), .ZN(n90) );
  OAI22_X1 U63 ( .A1(n38), .A2(n80), .B1(net108197), .B2(n36), .ZN(n31) );
  INV_X1 U64 ( .A(data_in[3]), .ZN(n80) );
  OAI22_X1 U65 ( .A1(n39), .A2(n70), .B1(net108198), .B2(n36), .ZN(n30) );
  INV_X1 U66 ( .A(data_in[4]), .ZN(n70) );
  OAI22_X1 U67 ( .A1(n39), .A2(n67), .B1(net108199), .B2(n36), .ZN(n29) );
  INV_X1 U68 ( .A(data_in[5]), .ZN(n67) );
  OAI22_X1 U69 ( .A1(n39), .A2(n66), .B1(net108200), .B2(n36), .ZN(n28) );
  INV_X1 U70 ( .A(data_in[6]), .ZN(n66) );
  OAI22_X1 U71 ( .A1(n39), .A2(n65), .B1(net108201), .B2(n36), .ZN(n27) );
  INV_X1 U72 ( .A(data_in[7]), .ZN(n65) );
  OAI22_X1 U73 ( .A1(n39), .A2(n64), .B1(net108202), .B2(n36), .ZN(n26) );
  INV_X1 U74 ( .A(data_in[8]), .ZN(n64) );
  OAI22_X1 U75 ( .A1(n40), .A2(n63), .B1(net108203), .B2(n36), .ZN(n25) );
  INV_X1 U76 ( .A(data_in[9]), .ZN(n63) );
  OAI22_X1 U77 ( .A1(n40), .A2(n62), .B1(net108204), .B2(n36), .ZN(n24) );
  INV_X1 U78 ( .A(data_in[10]), .ZN(n62) );
  OAI22_X1 U79 ( .A1(n40), .A2(n61), .B1(net108205), .B2(n36), .ZN(n23) );
  INV_X1 U80 ( .A(data_in[11]), .ZN(n61) );
endmodule


module NRegister_N32_39 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108194, net108195, net108196, net108197, net108198,
         net108199, net108200, net108201, net108202, net108203, net108204,
         net108205, net108206, net108207, net108208, net108209, net108210,
         net108211, net108212, net108213, net108214, net108215, net108216,
         net108217, net108218, net108219, net108220, net108221, net108222,
         net108223, net108224, net108225, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n46), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n46), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n46), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n44), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n46), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n44), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n44), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n44), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n46), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n44), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n44), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n44), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n44), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n44), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n44), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n44), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n44), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n45), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n45), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n45), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n45), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n45), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n45), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n45), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n45), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n45), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n46), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n46), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n46), .Q(data_out[0]), 
        .QN(net108194) );
  BUF_X1 U3 ( .A(n47), .Z(n45) );
  BUF_X1 U4 ( .A(n47), .Z(n44) );
  BUF_X1 U5 ( .A(n47), .Z(n46) );
  INV_X1 U6 ( .A(reset), .ZN(n47) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n92), .Z(n39) );
  BUF_X1 U10 ( .A(n92), .Z(n40) );
  BUF_X1 U11 ( .A(n92), .Z(n42) );
  BUF_X1 U12 ( .A(n92), .Z(n37) );
  BUF_X1 U13 ( .A(n92), .Z(n38) );
  BUF_X1 U14 ( .A(n92), .Z(n41) );
  BUF_X1 U15 ( .A(n92), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n85), .B1(net108194), .B2(n36), .ZN(n34) );
  INV_X1 U17 ( .A(data_in[0]), .ZN(n85) );
  OAI22_X1 U18 ( .A1(n38), .A2(n86), .B1(net108224), .B2(n35), .ZN(n4) );
  INV_X1 U19 ( .A(data_in[30]), .ZN(n86) );
  OAI22_X1 U20 ( .A1(n38), .A2(n83), .B1(net108196), .B2(n36), .ZN(n32) );
  INV_X1 U21 ( .A(data_in[2]), .ZN(n83) );
  OAI22_X1 U22 ( .A1(n38), .A2(n82), .B1(net108197), .B2(n36), .ZN(n31) );
  INV_X1 U23 ( .A(data_in[3]), .ZN(n82) );
  OAI22_X1 U24 ( .A1(n39), .A2(n81), .B1(net108198), .B2(n36), .ZN(n30) );
  INV_X1 U25 ( .A(data_in[4]), .ZN(n81) );
  OAI22_X1 U26 ( .A1(n39), .A2(n70), .B1(net108199), .B2(n36), .ZN(n29) );
  INV_X1 U27 ( .A(data_in[5]), .ZN(n70) );
  OAI22_X1 U28 ( .A1(n39), .A2(n67), .B1(net108200), .B2(n36), .ZN(n28) );
  INV_X1 U29 ( .A(data_in[6]), .ZN(n67) );
  OAI22_X1 U30 ( .A1(n39), .A2(n66), .B1(net108201), .B2(n36), .ZN(n27) );
  INV_X1 U31 ( .A(data_in[7]), .ZN(n66) );
  OAI22_X1 U32 ( .A1(n41), .A2(n58), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U33 ( .A(data_in[31]), .ZN(n58) );
  OAI22_X1 U34 ( .A1(n38), .A2(n84), .B1(net108195), .B2(n36), .ZN(n33) );
  INV_X1 U35 ( .A(data_in[1]), .ZN(n84) );
  OAI22_X1 U36 ( .A1(n39), .A2(n65), .B1(net108202), .B2(n36), .ZN(n26) );
  INV_X1 U37 ( .A(data_in[8]), .ZN(n65) );
  OAI22_X1 U38 ( .A1(n40), .A2(n64), .B1(net108203), .B2(n36), .ZN(n25) );
  INV_X1 U39 ( .A(data_in[9]), .ZN(n64) );
  OAI22_X1 U40 ( .A1(n40), .A2(n63), .B1(net108204), .B2(n36), .ZN(n24) );
  INV_X1 U41 ( .A(data_in[10]), .ZN(n63) );
  OAI22_X1 U42 ( .A1(n40), .A2(n62), .B1(net108205), .B2(n36), .ZN(n23) );
  INV_X1 U43 ( .A(data_in[11]), .ZN(n62) );
  OAI22_X1 U44 ( .A1(n40), .A2(n61), .B1(net108206), .B2(n36), .ZN(n22) );
  INV_X1 U45 ( .A(data_in[12]), .ZN(n61) );
  OAI22_X1 U46 ( .A1(n40), .A2(n60), .B1(net108207), .B2(n36), .ZN(n21) );
  INV_X1 U47 ( .A(data_in[13]), .ZN(n60) );
  OAI22_X1 U48 ( .A1(n41), .A2(n59), .B1(net108208), .B2(n35), .ZN(n20) );
  INV_X1 U49 ( .A(data_in[14]), .ZN(n59) );
  OAI22_X1 U50 ( .A1(n41), .A2(n57), .B1(net108209), .B2(n35), .ZN(n19) );
  INV_X1 U51 ( .A(data_in[15]), .ZN(n57) );
  OAI22_X1 U52 ( .A1(n41), .A2(n56), .B1(net108210), .B2(n35), .ZN(n18) );
  INV_X1 U53 ( .A(data_in[16]), .ZN(n56) );
  OAI22_X1 U54 ( .A1(n41), .A2(n55), .B1(net108211), .B2(n35), .ZN(n17) );
  INV_X1 U55 ( .A(data_in[17]), .ZN(n55) );
  OAI22_X1 U56 ( .A1(n42), .A2(n54), .B1(net108212), .B2(n35), .ZN(n16) );
  INV_X1 U57 ( .A(data_in[18]), .ZN(n54) );
  OAI22_X1 U58 ( .A1(n42), .A2(n53), .B1(net108213), .B2(n35), .ZN(n15) );
  INV_X1 U59 ( .A(data_in[19]), .ZN(n53) );
  OAI22_X1 U60 ( .A1(n42), .A2(n52), .B1(net108214), .B2(n35), .ZN(n14) );
  INV_X1 U61 ( .A(data_in[20]), .ZN(n52) );
  OAI22_X1 U62 ( .A1(n42), .A2(n51), .B1(net108215), .B2(n35), .ZN(n13) );
  INV_X1 U63 ( .A(data_in[21]), .ZN(n51) );
  OAI22_X1 U64 ( .A1(n42), .A2(n50), .B1(net108216), .B2(n35), .ZN(n12) );
  INV_X1 U65 ( .A(data_in[22]), .ZN(n50) );
  OAI22_X1 U66 ( .A1(n43), .A2(n49), .B1(net108217), .B2(n35), .ZN(n11) );
  INV_X1 U67 ( .A(data_in[23]), .ZN(n49) );
  OAI22_X1 U68 ( .A1(n43), .A2(n48), .B1(net108218), .B2(n35), .ZN(n10) );
  INV_X1 U69 ( .A(data_in[24]), .ZN(n48) );
  OAI22_X1 U70 ( .A1(n37), .A2(n91), .B1(net108219), .B2(n35), .ZN(n9) );
  INV_X1 U71 ( .A(data_in[25]), .ZN(n91) );
  OAI22_X1 U72 ( .A1(n37), .A2(n90), .B1(net108220), .B2(n36), .ZN(n8) );
  INV_X1 U73 ( .A(data_in[26]), .ZN(n90) );
  OAI22_X1 U74 ( .A1(n37), .A2(n89), .B1(net108221), .B2(n35), .ZN(n7) );
  INV_X1 U75 ( .A(data_in[27]), .ZN(n89) );
  OAI22_X1 U76 ( .A1(n37), .A2(n88), .B1(net108222), .B2(n36), .ZN(n6) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n88) );
  OAI22_X1 U78 ( .A1(n37), .A2(n87), .B1(net108223), .B2(n35), .ZN(n5) );
  INV_X1 U79 ( .A(data_in[29]), .ZN(n87) );
  NAND2_X1 U80 ( .A1(load), .A2(enable), .ZN(n92) );
endmodule


module NRegister_N32_38 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108194, net108195, net108196, net108197, net108198,
         net108199, net108200, net108201, net108202, net108203, net108204,
         net108205, net108206, net108207, net108208, net108209, net108210,
         net108211, net108212, net108213, net108214, net108215, net108216,
         net108217, net108218, net108219, net108220, net108221, net108222,
         net108223, net108224, net108225, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n46), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n46), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n46), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n44), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n46), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n44), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n44), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n44), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n46), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n44), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n44), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n44), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n44), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n44), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n44), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n44), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n44), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n45), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n45), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n45), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n45), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n45), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n45), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n45), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n45), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n45), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n46), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n46), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n46), .Q(data_out[0]), 
        .QN(net108194) );
  BUF_X1 U3 ( .A(n47), .Z(n45) );
  BUF_X1 U4 ( .A(n47), .Z(n44) );
  BUF_X1 U5 ( .A(n47), .Z(n46) );
  INV_X1 U6 ( .A(reset), .ZN(n47) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n92), .Z(n39) );
  BUF_X1 U10 ( .A(n92), .Z(n40) );
  BUF_X1 U11 ( .A(n92), .Z(n42) );
  BUF_X1 U12 ( .A(n92), .Z(n37) );
  BUF_X1 U13 ( .A(n92), .Z(n38) );
  BUF_X1 U14 ( .A(n92), .Z(n41) );
  BUF_X1 U15 ( .A(n92), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n85), .B1(net108194), .B2(n36), .ZN(n34) );
  INV_X1 U17 ( .A(data_in[0]), .ZN(n85) );
  OAI22_X1 U18 ( .A1(n38), .A2(n84), .B1(net108195), .B2(n35), .ZN(n33) );
  INV_X1 U19 ( .A(data_in[1]), .ZN(n84) );
  OAI22_X1 U20 ( .A1(n37), .A2(n91), .B1(net108219), .B2(n36), .ZN(n9) );
  INV_X1 U21 ( .A(data_in[25]), .ZN(n91) );
  OAI22_X1 U22 ( .A1(n37), .A2(n90), .B1(net108220), .B2(n35), .ZN(n8) );
  INV_X1 U23 ( .A(data_in[26]), .ZN(n90) );
  OAI22_X1 U24 ( .A1(n37), .A2(n89), .B1(net108221), .B2(n36), .ZN(n7) );
  INV_X1 U25 ( .A(data_in[27]), .ZN(n89) );
  OAI22_X1 U26 ( .A1(n37), .A2(n88), .B1(net108222), .B2(n35), .ZN(n6) );
  INV_X1 U27 ( .A(data_in[28]), .ZN(n88) );
  OAI22_X1 U28 ( .A1(n37), .A2(n87), .B1(net108223), .B2(n36), .ZN(n5) );
  INV_X1 U29 ( .A(data_in[29]), .ZN(n87) );
  OAI22_X1 U30 ( .A1(n38), .A2(n86), .B1(net108224), .B2(n35), .ZN(n4) );
  INV_X1 U31 ( .A(data_in[30]), .ZN(n86) );
  OAI22_X1 U32 ( .A1(n38), .A2(n83), .B1(net108196), .B2(n36), .ZN(n32) );
  INV_X1 U33 ( .A(data_in[2]), .ZN(n83) );
  OAI22_X1 U34 ( .A1(n38), .A2(n82), .B1(net108197), .B2(n36), .ZN(n31) );
  INV_X1 U35 ( .A(data_in[3]), .ZN(n82) );
  OAI22_X1 U36 ( .A1(n39), .A2(n81), .B1(net108198), .B2(n36), .ZN(n30) );
  INV_X1 U37 ( .A(data_in[4]), .ZN(n81) );
  OAI22_X1 U38 ( .A1(n39), .A2(n70), .B1(net108199), .B2(n36), .ZN(n29) );
  INV_X1 U39 ( .A(data_in[5]), .ZN(n70) );
  OAI22_X1 U40 ( .A1(n39), .A2(n67), .B1(net108200), .B2(n36), .ZN(n28) );
  INV_X1 U41 ( .A(data_in[6]), .ZN(n67) );
  OAI22_X1 U42 ( .A1(n39), .A2(n66), .B1(net108201), .B2(n36), .ZN(n27) );
  INV_X1 U43 ( .A(data_in[7]), .ZN(n66) );
  OAI22_X1 U44 ( .A1(n39), .A2(n65), .B1(net108202), .B2(n36), .ZN(n26) );
  INV_X1 U45 ( .A(data_in[8]), .ZN(n65) );
  OAI22_X1 U46 ( .A1(n40), .A2(n64), .B1(net108203), .B2(n36), .ZN(n25) );
  INV_X1 U47 ( .A(data_in[9]), .ZN(n64) );
  OAI22_X1 U48 ( .A1(n40), .A2(n63), .B1(net108204), .B2(n36), .ZN(n24) );
  INV_X1 U49 ( .A(data_in[10]), .ZN(n63) );
  OAI22_X1 U50 ( .A1(n40), .A2(n62), .B1(net108205), .B2(n36), .ZN(n23) );
  INV_X1 U51 ( .A(data_in[11]), .ZN(n62) );
  OAI22_X1 U52 ( .A1(n40), .A2(n61), .B1(net108206), .B2(n36), .ZN(n22) );
  INV_X1 U53 ( .A(data_in[12]), .ZN(n61) );
  OAI22_X1 U54 ( .A1(n40), .A2(n60), .B1(net108207), .B2(n36), .ZN(n21) );
  INV_X1 U55 ( .A(data_in[13]), .ZN(n60) );
  OAI22_X1 U56 ( .A1(n41), .A2(n59), .B1(net108208), .B2(n35), .ZN(n20) );
  INV_X1 U57 ( .A(data_in[14]), .ZN(n59) );
  OAI22_X1 U58 ( .A1(n41), .A2(n57), .B1(net108209), .B2(n35), .ZN(n19) );
  INV_X1 U59 ( .A(data_in[15]), .ZN(n57) );
  OAI22_X1 U60 ( .A1(n41), .A2(n56), .B1(net108210), .B2(n35), .ZN(n18) );
  INV_X1 U61 ( .A(data_in[16]), .ZN(n56) );
  OAI22_X1 U62 ( .A1(n41), .A2(n55), .B1(net108211), .B2(n35), .ZN(n17) );
  INV_X1 U63 ( .A(data_in[17]), .ZN(n55) );
  OAI22_X1 U64 ( .A1(n42), .A2(n54), .B1(net108212), .B2(n35), .ZN(n16) );
  INV_X1 U65 ( .A(data_in[18]), .ZN(n54) );
  OAI22_X1 U66 ( .A1(n42), .A2(n53), .B1(net108213), .B2(n35), .ZN(n15) );
  INV_X1 U67 ( .A(data_in[19]), .ZN(n53) );
  OAI22_X1 U68 ( .A1(n42), .A2(n52), .B1(net108214), .B2(n35), .ZN(n14) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n52) );
  OAI22_X1 U70 ( .A1(n42), .A2(n51), .B1(net108215), .B2(n35), .ZN(n13) );
  INV_X1 U71 ( .A(data_in[21]), .ZN(n51) );
  OAI22_X1 U72 ( .A1(n42), .A2(n50), .B1(net108216), .B2(n35), .ZN(n12) );
  INV_X1 U73 ( .A(data_in[22]), .ZN(n50) );
  OAI22_X1 U74 ( .A1(n43), .A2(n49), .B1(net108217), .B2(n35), .ZN(n11) );
  INV_X1 U75 ( .A(data_in[23]), .ZN(n49) );
  OAI22_X1 U76 ( .A1(n43), .A2(n48), .B1(net108218), .B2(n35), .ZN(n10) );
  INV_X1 U77 ( .A(data_in[24]), .ZN(n48) );
  OAI22_X1 U78 ( .A1(n41), .A2(n58), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U79 ( .A(data_in[31]), .ZN(n58) );
  NAND2_X1 U80 ( .A1(load), .A2(enable), .ZN(n92) );
endmodule


module NRegister_N32_37 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108194, net108195, net108196, net108197, net108198,
         net108199, net108200, net108201, net108202, net108203, net108204,
         net108205, net108206, net108207, net108208, net108209, net108210,
         net108211, net108212, net108213, net108214, net108215, net108216,
         net108217, net108218, net108219, net108220, net108221, net108222,
         net108223, net108224, net108225, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n46), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n46), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n46), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n44), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n46), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n44), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n44), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n44), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n46), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n44), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n44), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n44), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n44), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n44), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n44), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n44), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n44), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n45), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n45), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n45), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n45), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n45), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n45), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n45), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n45), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n45), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n46), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n46), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n46), .Q(data_out[0]), 
        .QN(net108194) );
  BUF_X1 U3 ( .A(n47), .Z(n45) );
  BUF_X1 U4 ( .A(n47), .Z(n44) );
  BUF_X1 U5 ( .A(n47), .Z(n46) );
  INV_X1 U6 ( .A(reset), .ZN(n47) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n92), .Z(n39) );
  BUF_X1 U10 ( .A(n92), .Z(n40) );
  BUF_X1 U11 ( .A(n92), .Z(n42) );
  BUF_X1 U12 ( .A(n92), .Z(n37) );
  BUF_X1 U13 ( .A(n92), .Z(n38) );
  BUF_X1 U14 ( .A(n92), .Z(n41) );
  BUF_X1 U15 ( .A(n92), .Z(n43) );
  OAI22_X1 U16 ( .A1(n38), .A2(n85), .B1(net108194), .B2(n36), .ZN(n34) );
  INV_X1 U17 ( .A(data_in[0]), .ZN(n85) );
  OAI22_X1 U18 ( .A1(n38), .A2(n84), .B1(net108195), .B2(n35), .ZN(n33) );
  INV_X1 U19 ( .A(data_in[1]), .ZN(n84) );
  OAI22_X1 U20 ( .A1(n37), .A2(n91), .B1(net108219), .B2(n36), .ZN(n9) );
  INV_X1 U21 ( .A(data_in[25]), .ZN(n91) );
  OAI22_X1 U22 ( .A1(n38), .A2(n83), .B1(net108196), .B2(n36), .ZN(n32) );
  INV_X1 U23 ( .A(data_in[2]), .ZN(n83) );
  OAI22_X1 U24 ( .A1(n38), .A2(n82), .B1(net108197), .B2(n36), .ZN(n31) );
  INV_X1 U25 ( .A(data_in[3]), .ZN(n82) );
  OAI22_X1 U26 ( .A1(n39), .A2(n81), .B1(net108198), .B2(n36), .ZN(n30) );
  INV_X1 U27 ( .A(data_in[4]), .ZN(n81) );
  OAI22_X1 U28 ( .A1(n39), .A2(n70), .B1(net108199), .B2(n36), .ZN(n29) );
  INV_X1 U29 ( .A(data_in[5]), .ZN(n70) );
  OAI22_X1 U30 ( .A1(n39), .A2(n67), .B1(net108200), .B2(n36), .ZN(n28) );
  INV_X1 U31 ( .A(data_in[6]), .ZN(n67) );
  OAI22_X1 U32 ( .A1(n39), .A2(n66), .B1(net108201), .B2(n36), .ZN(n27) );
  INV_X1 U33 ( .A(data_in[7]), .ZN(n66) );
  OAI22_X1 U34 ( .A1(n39), .A2(n65), .B1(net108202), .B2(n36), .ZN(n26) );
  INV_X1 U35 ( .A(data_in[8]), .ZN(n65) );
  OAI22_X1 U36 ( .A1(n40), .A2(n64), .B1(net108203), .B2(n36), .ZN(n25) );
  INV_X1 U37 ( .A(data_in[9]), .ZN(n64) );
  OAI22_X1 U38 ( .A1(n40), .A2(n63), .B1(net108204), .B2(n36), .ZN(n24) );
  INV_X1 U39 ( .A(data_in[10]), .ZN(n63) );
  OAI22_X1 U40 ( .A1(n40), .A2(n62), .B1(net108205), .B2(n36), .ZN(n23) );
  INV_X1 U41 ( .A(data_in[11]), .ZN(n62) );
  OAI22_X1 U42 ( .A1(n40), .A2(n61), .B1(net108206), .B2(n36), .ZN(n22) );
  INV_X1 U43 ( .A(data_in[12]), .ZN(n61) );
  OAI22_X1 U44 ( .A1(n40), .A2(n60), .B1(net108207), .B2(n36), .ZN(n21) );
  INV_X1 U45 ( .A(data_in[13]), .ZN(n60) );
  OAI22_X1 U46 ( .A1(n41), .A2(n59), .B1(net108208), .B2(n35), .ZN(n20) );
  INV_X1 U47 ( .A(data_in[14]), .ZN(n59) );
  OAI22_X1 U48 ( .A1(n41), .A2(n57), .B1(net108209), .B2(n35), .ZN(n19) );
  INV_X1 U49 ( .A(data_in[15]), .ZN(n57) );
  OAI22_X1 U50 ( .A1(n43), .A2(n49), .B1(net108217), .B2(n35), .ZN(n11) );
  INV_X1 U51 ( .A(data_in[23]), .ZN(n49) );
  NAND2_X1 U52 ( .A1(load), .A2(enable), .ZN(n92) );
  OAI22_X1 U53 ( .A1(n42), .A2(n52), .B1(net108214), .B2(n35), .ZN(n14) );
  INV_X1 U54 ( .A(data_in[20]), .ZN(n52) );
  OAI22_X1 U55 ( .A1(n42), .A2(n51), .B1(net108215), .B2(n35), .ZN(n13) );
  INV_X1 U56 ( .A(data_in[21]), .ZN(n51) );
  OAI22_X1 U57 ( .A1(n42), .A2(n50), .B1(net108216), .B2(n35), .ZN(n12) );
  INV_X1 U58 ( .A(data_in[22]), .ZN(n50) );
  OAI22_X1 U59 ( .A1(n43), .A2(n48), .B1(net108218), .B2(n35), .ZN(n10) );
  INV_X1 U60 ( .A(data_in[24]), .ZN(n48) );
  OAI22_X1 U61 ( .A1(n41), .A2(n56), .B1(net108210), .B2(n35), .ZN(n18) );
  INV_X1 U62 ( .A(data_in[16]), .ZN(n56) );
  OAI22_X1 U63 ( .A1(n41), .A2(n55), .B1(net108211), .B2(n35), .ZN(n17) );
  INV_X1 U64 ( .A(data_in[17]), .ZN(n55) );
  OAI22_X1 U65 ( .A1(n42), .A2(n54), .B1(net108212), .B2(n35), .ZN(n16) );
  INV_X1 U66 ( .A(data_in[18]), .ZN(n54) );
  OAI22_X1 U67 ( .A1(n42), .A2(n53), .B1(net108213), .B2(n35), .ZN(n15) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n53) );
  OAI22_X1 U69 ( .A1(n37), .A2(n90), .B1(net108220), .B2(n35), .ZN(n8) );
  INV_X1 U70 ( .A(data_in[26]), .ZN(n90) );
  OAI22_X1 U71 ( .A1(n37), .A2(n89), .B1(net108221), .B2(n36), .ZN(n7) );
  INV_X1 U72 ( .A(data_in[27]), .ZN(n89) );
  OAI22_X1 U73 ( .A1(n37), .A2(n88), .B1(net108222), .B2(n35), .ZN(n6) );
  INV_X1 U74 ( .A(data_in[28]), .ZN(n88) );
  OAI22_X1 U75 ( .A1(n37), .A2(n87), .B1(net108223), .B2(n36), .ZN(n5) );
  INV_X1 U76 ( .A(data_in[29]), .ZN(n87) );
  OAI22_X1 U77 ( .A1(n38), .A2(n86), .B1(net108224), .B2(n35), .ZN(n4) );
  INV_X1 U78 ( .A(data_in[30]), .ZN(n86) );
  OAI22_X1 U79 ( .A1(n41), .A2(n58), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n58) );
endmodule


module NRegister_N32_36 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, net108194, net108195, net108196, net108197,
         net108198, net108199, net108200, net108201, net108202, net108203,
         net108204, net108205, net108206, net108207, net108208, net108209,
         net108210, net108211, net108212, net108213, net108214, net108215,
         net108216, net108217, net108218, net108219, net108220, net108221,
         net108222, net108223, net108224, net108225, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n70, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n44), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n44), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n44), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n46), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n44), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n46), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n46), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n46), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n44), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n46), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n46), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n46), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n46), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n45), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n45), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n45), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n45), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n45), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n45), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n45), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n45), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n45), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n44), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n44), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n44), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n44), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n44), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n44), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n44), .Q(data_out[0]), 
        .QN(net108194) );
  INV_X1 U3 ( .A(n43), .ZN(n36) );
  INV_X1 U4 ( .A(n43), .ZN(n35) );
  BUF_X1 U5 ( .A(n90), .Z(n39) );
  BUF_X1 U6 ( .A(n90), .Z(n40) );
  BUF_X1 U7 ( .A(n90), .Z(n42) );
  BUF_X1 U8 ( .A(n90), .Z(n37) );
  BUF_X1 U9 ( .A(n90), .Z(n38) );
  BUF_X1 U10 ( .A(n90), .Z(n41) );
  BUF_X1 U11 ( .A(n90), .Z(n43) );
  BUF_X1 U12 ( .A(n3), .Z(n45) );
  BUF_X1 U13 ( .A(n3), .Z(n44) );
  BUF_X1 U14 ( .A(n3), .Z(n46) );
  OAI22_X1 U15 ( .A1(n37), .A2(n85), .B1(net108223), .B2(n36), .ZN(n5) );
  INV_X1 U16 ( .A(data_in[29]), .ZN(n85) );
  OAI22_X1 U17 ( .A1(n38), .A2(n84), .B1(net108224), .B2(n35), .ZN(n4) );
  INV_X1 U18 ( .A(data_in[30]), .ZN(n84) );
  OAI22_X1 U19 ( .A1(n37), .A2(n89), .B1(net108219), .B2(n36), .ZN(n9) );
  INV_X1 U20 ( .A(data_in[25]), .ZN(n89) );
  OAI22_X1 U21 ( .A1(n37), .A2(n88), .B1(net108220), .B2(n35), .ZN(n8) );
  INV_X1 U22 ( .A(data_in[26]), .ZN(n88) );
  OAI22_X1 U23 ( .A1(n37), .A2(n87), .B1(net108221), .B2(n36), .ZN(n7) );
  INV_X1 U24 ( .A(data_in[27]), .ZN(n87) );
  OAI22_X1 U25 ( .A1(n37), .A2(n86), .B1(net108222), .B2(n35), .ZN(n6) );
  INV_X1 U26 ( .A(data_in[28]), .ZN(n86) );
  OAI22_X1 U27 ( .A1(n41), .A2(n57), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U28 ( .A(data_in[31]), .ZN(n57) );
  OAI22_X1 U29 ( .A1(n43), .A2(n48), .B1(net108217), .B2(n35), .ZN(n11) );
  INV_X1 U30 ( .A(data_in[23]), .ZN(n48) );
  OAI22_X1 U31 ( .A1(n43), .A2(n47), .B1(net108218), .B2(n35), .ZN(n10) );
  INV_X1 U32 ( .A(data_in[24]), .ZN(n47) );
  OAI22_X1 U33 ( .A1(n42), .A2(n49), .B1(net108216), .B2(n35), .ZN(n12) );
  INV_X1 U34 ( .A(data_in[22]), .ZN(n49) );
  OAI22_X1 U35 ( .A1(n41), .A2(n58), .B1(net108208), .B2(n35), .ZN(n20) );
  INV_X1 U36 ( .A(data_in[14]), .ZN(n58) );
  OAI22_X1 U37 ( .A1(n41), .A2(n56), .B1(net108209), .B2(n35), .ZN(n19) );
  INV_X1 U38 ( .A(data_in[15]), .ZN(n56) );
  OAI22_X1 U39 ( .A1(n41), .A2(n54), .B1(net108211), .B2(n35), .ZN(n17) );
  INV_X1 U40 ( .A(data_in[17]), .ZN(n54) );
  OAI22_X1 U41 ( .A1(n42), .A2(n52), .B1(net108213), .B2(n35), .ZN(n15) );
  INV_X1 U42 ( .A(data_in[19]), .ZN(n52) );
  OAI22_X1 U43 ( .A1(n42), .A2(n50), .B1(net108215), .B2(n35), .ZN(n13) );
  INV_X1 U44 ( .A(data_in[21]), .ZN(n50) );
  OAI22_X1 U45 ( .A1(n41), .A2(n55), .B1(net108210), .B2(n35), .ZN(n18) );
  INV_X1 U46 ( .A(data_in[16]), .ZN(n55) );
  OAI22_X1 U47 ( .A1(n42), .A2(n53), .B1(net108212), .B2(n35), .ZN(n16) );
  INV_X1 U48 ( .A(data_in[18]), .ZN(n53) );
  OAI22_X1 U49 ( .A1(n42), .A2(n51), .B1(net108214), .B2(n35), .ZN(n14) );
  INV_X1 U50 ( .A(data_in[20]), .ZN(n51) );
  OAI22_X1 U51 ( .A1(n39), .A2(n65), .B1(net108201), .B2(n36), .ZN(n27) );
  INV_X1 U52 ( .A(data_in[7]), .ZN(n65) );
  OAI22_X1 U53 ( .A1(n40), .A2(n63), .B1(net108203), .B2(n36), .ZN(n25) );
  INV_X1 U54 ( .A(data_in[9]), .ZN(n63) );
  OAI22_X1 U55 ( .A1(n40), .A2(n62), .B1(net108204), .B2(n36), .ZN(n24) );
  INV_X1 U56 ( .A(data_in[10]), .ZN(n62) );
  OAI22_X1 U57 ( .A1(n40), .A2(n61), .B1(net108205), .B2(n36), .ZN(n23) );
  INV_X1 U58 ( .A(data_in[11]), .ZN(n61) );
  OAI22_X1 U59 ( .A1(n40), .A2(n59), .B1(net108207), .B2(n36), .ZN(n21) );
  INV_X1 U60 ( .A(data_in[13]), .ZN(n59) );
  OAI22_X1 U61 ( .A1(n39), .A2(n66), .B1(net108200), .B2(n36), .ZN(n28) );
  INV_X1 U62 ( .A(data_in[6]), .ZN(n66) );
  OAI22_X1 U63 ( .A1(n39), .A2(n64), .B1(net108202), .B2(n36), .ZN(n26) );
  INV_X1 U64 ( .A(data_in[8]), .ZN(n64) );
  OAI22_X1 U65 ( .A1(n40), .A2(n60), .B1(net108206), .B2(n36), .ZN(n22) );
  INV_X1 U66 ( .A(data_in[12]), .ZN(n60) );
  OAI22_X1 U67 ( .A1(n38), .A2(n81), .B1(net108196), .B2(n36), .ZN(n32) );
  INV_X1 U68 ( .A(data_in[2]), .ZN(n81) );
  OAI22_X1 U69 ( .A1(n38), .A2(n80), .B1(net108197), .B2(n36), .ZN(n31) );
  INV_X1 U70 ( .A(data_in[3]), .ZN(n80) );
  OAI22_X1 U71 ( .A1(n39), .A2(n70), .B1(net108198), .B2(n36), .ZN(n30) );
  INV_X1 U72 ( .A(data_in[4]), .ZN(n70) );
  OAI22_X1 U73 ( .A1(n38), .A2(n83), .B1(net108194), .B2(n36), .ZN(n34) );
  INV_X1 U74 ( .A(data_in[0]), .ZN(n83) );
  OAI22_X1 U75 ( .A1(n38), .A2(n82), .B1(net108195), .B2(n35), .ZN(n33) );
  INV_X1 U76 ( .A(data_in[1]), .ZN(n82) );
  OAI22_X1 U77 ( .A1(n39), .A2(n67), .B1(net108199), .B2(n36), .ZN(n29) );
  INV_X1 U78 ( .A(data_in[5]), .ZN(n67) );
  NAND2_X1 U79 ( .A1(load), .A2(enable), .ZN(n90) );
  INV_X1 U80 ( .A(reset), .ZN(n3) );
endmodule


module NRegister_N32_35 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108194, net108195, net108196, net108197, net108198,
         net108199, net108200, net108201, net108202, net108203, net108204,
         net108205, net108206, net108207, net108208, net108209, net108210,
         net108211, net108212, net108213, net108214, net108215, net108216,
         net108217, net108218, net108219, net108220, net108221, net108222,
         net108223, net108224, net108225, n68, net145577, net145575, net145573,
         net145571, net145569, net145567, net145565, net145563, net145561,
         net145559, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n70, n73, n74, n75;

  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n38), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n40), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n38), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n40), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n40), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n40), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n40), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n39), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n39), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n39), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n39), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n39), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n39), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n39), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n39), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n39), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n39), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n39), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n39), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n38), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n38), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n38), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n38), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n38), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n38), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n38), .Q(data_out[0]), 
        .QN(net108194) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n40), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n40), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X2 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n38), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X2 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n38), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X2 \data_out_reg[31]  ( .D(n35), .CK(clk), .RN(n38), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X2 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n40), .Q(data_out[25]), 
        .QN(net108219) );
  BUF_X1 U3 ( .A(n68), .Z(net145567) );
  INV_X1 U4 ( .A(net145577), .ZN(net145559) );
  BUF_X1 U5 ( .A(n68), .Z(net145565) );
  OR2_X1 U6 ( .A1(net108225), .A2(net145559), .ZN(n36) );
  BUF_X1 U7 ( .A(n68), .Z(net145573) );
  INV_X1 U8 ( .A(net145577), .ZN(net145563) );
  NAND2_X1 U9 ( .A1(n37), .A2(n36), .ZN(n35) );
  NAND2_X1 U10 ( .A1(data_in[31]), .A2(net145563), .ZN(n37) );
  BUF_X1 U11 ( .A(n68), .Z(net145577) );
  NAND2_X1 U12 ( .A1(load), .A2(enable), .ZN(n68) );
  INV_X1 U13 ( .A(net145577), .ZN(net145561) );
  BUF_X1 U14 ( .A(n68), .Z(net145569) );
  BUF_X1 U15 ( .A(n68), .Z(net145571) );
  BUF_X1 U16 ( .A(n68), .Z(net145575) );
  BUF_X1 U17 ( .A(n3), .Z(n39) );
  BUF_X1 U18 ( .A(n3), .Z(n38) );
  BUF_X1 U19 ( .A(n3), .Z(n40) );
  OAI22_X1 U20 ( .A1(n66), .A2(net145567), .B1(net108224), .B2(net145563), 
        .ZN(n4) );
  INV_X1 U21 ( .A(data_in[30]), .ZN(n66) );
  OAI22_X1 U22 ( .A1(n67), .A2(net145565), .B1(net108223), .B2(net145563), 
        .ZN(n5) );
  INV_X1 U23 ( .A(data_in[29]), .ZN(n67) );
  OAI22_X1 U24 ( .A1(n70), .A2(net145565), .B1(net108222), .B2(net145563), 
        .ZN(n6) );
  INV_X1 U25 ( .A(data_in[28]), .ZN(n70) );
  OAI22_X1 U26 ( .A1(n73), .A2(net145565), .B1(net108221), .B2(net145563), 
        .ZN(n7) );
  INV_X1 U27 ( .A(data_in[27]), .ZN(n73) );
  OAI22_X1 U28 ( .A1(n74), .A2(net145565), .B1(net108220), .B2(net145563), 
        .ZN(n8) );
  INV_X1 U29 ( .A(data_in[26]), .ZN(n74) );
  OAI22_X1 U30 ( .A1(n75), .A2(net145565), .B1(net108219), .B2(net145563), 
        .ZN(n9) );
  INV_X1 U31 ( .A(data_in[25]), .ZN(n75) );
  OAI22_X1 U32 ( .A1(n41), .A2(net145577), .B1(net108218), .B2(net145559), 
        .ZN(n10) );
  INV_X1 U33 ( .A(data_in[24]), .ZN(n41) );
  OAI22_X1 U34 ( .A1(net145577), .A2(n42), .B1(net108217), .B2(net145559), 
        .ZN(n11) );
  INV_X1 U35 ( .A(data_in[23]), .ZN(n42) );
  OAI22_X1 U36 ( .A1(net145575), .A2(n43), .B1(net108216), .B2(net145559), 
        .ZN(n12) );
  INV_X1 U37 ( .A(data_in[22]), .ZN(n43) );
  OAI22_X1 U38 ( .A1(net145575), .A2(n44), .B1(net108215), .B2(net145559), 
        .ZN(n13) );
  INV_X1 U39 ( .A(data_in[21]), .ZN(n44) );
  OAI22_X1 U40 ( .A1(net145567), .A2(n64), .B1(net108195), .B2(net145563), 
        .ZN(n33) );
  INV_X1 U41 ( .A(data_in[1]), .ZN(n64) );
  OAI22_X1 U42 ( .A1(net145567), .A2(n65), .B1(net108194), .B2(net145563), 
        .ZN(n34) );
  INV_X1 U43 ( .A(data_in[0]), .ZN(n65) );
  OAI22_X1 U44 ( .A1(net145569), .A2(n59), .B1(net108200), .B2(net145561), 
        .ZN(n28) );
  INV_X1 U45 ( .A(data_in[6]), .ZN(n59) );
  OAI22_X1 U46 ( .A1(net145571), .A2(n52), .B1(net108207), .B2(net145561), 
        .ZN(n21) );
  INV_X1 U47 ( .A(data_in[13]), .ZN(n52) );
  OAI22_X1 U48 ( .A1(net145571), .A2(n53), .B1(net108206), .B2(net145561), 
        .ZN(n22) );
  INV_X1 U49 ( .A(data_in[12]), .ZN(n53) );
  OAI22_X1 U50 ( .A1(net145571), .A2(n56), .B1(net108203), .B2(net145561), 
        .ZN(n25) );
  INV_X1 U51 ( .A(data_in[9]), .ZN(n56) );
  OAI22_X1 U52 ( .A1(net145571), .A2(n54), .B1(net108205), .B2(net145561), 
        .ZN(n23) );
  INV_X1 U53 ( .A(data_in[11]), .ZN(n54) );
  OAI22_X1 U54 ( .A1(net145569), .A2(n57), .B1(net108202), .B2(net145561), 
        .ZN(n26) );
  INV_X1 U55 ( .A(data_in[8]), .ZN(n57) );
  OAI22_X1 U56 ( .A1(net145571), .A2(n55), .B1(net108204), .B2(net145561), 
        .ZN(n24) );
  INV_X1 U57 ( .A(data_in[10]), .ZN(n55) );
  OAI22_X1 U58 ( .A1(net145569), .A2(n58), .B1(net108201), .B2(net145561), 
        .ZN(n27) );
  INV_X1 U59 ( .A(data_in[7]), .ZN(n58) );
  OAI22_X1 U60 ( .A1(net145569), .A2(n60), .B1(net108199), .B2(net145561), 
        .ZN(n29) );
  INV_X1 U61 ( .A(data_in[5]), .ZN(n60) );
  OAI22_X1 U62 ( .A1(net145569), .A2(n61), .B1(net108198), .B2(net145561), 
        .ZN(n30) );
  INV_X1 U63 ( .A(data_in[4]), .ZN(n61) );
  OAI22_X1 U64 ( .A1(net145567), .A2(n62), .B1(net108197), .B2(net145561), 
        .ZN(n31) );
  INV_X1 U65 ( .A(data_in[3]), .ZN(n62) );
  OAI22_X1 U66 ( .A1(net145567), .A2(n63), .B1(net108196), .B2(net145561), 
        .ZN(n32) );
  INV_X1 U67 ( .A(data_in[2]), .ZN(n63) );
  OAI22_X1 U68 ( .A1(net145575), .A2(n45), .B1(net108214), .B2(net145559), 
        .ZN(n14) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n45) );
  OAI22_X1 U70 ( .A1(net145575), .A2(n46), .B1(net108213), .B2(net145559), 
        .ZN(n15) );
  INV_X1 U71 ( .A(data_in[19]), .ZN(n46) );
  OAI22_X1 U72 ( .A1(net145573), .A2(n48), .B1(net108211), .B2(net145559), 
        .ZN(n17) );
  INV_X1 U73 ( .A(data_in[17]), .ZN(n48) );
  OAI22_X1 U74 ( .A1(net145575), .A2(n47), .B1(net108212), .B2(net145559), 
        .ZN(n16) );
  INV_X1 U75 ( .A(data_in[18]), .ZN(n47) );
  OAI22_X1 U76 ( .A1(net145573), .A2(n49), .B1(net108210), .B2(net145559), 
        .ZN(n18) );
  INV_X1 U77 ( .A(data_in[16]), .ZN(n49) );
  OAI22_X1 U78 ( .A1(net145573), .A2(n50), .B1(net108209), .B2(net145559), 
        .ZN(n19) );
  INV_X1 U79 ( .A(data_in[15]), .ZN(n50) );
  OAI22_X1 U80 ( .A1(net145573), .A2(n51), .B1(net108208), .B2(net145559), 
        .ZN(n20) );
  INV_X1 U81 ( .A(data_in[14]), .ZN(n51) );
  INV_X1 U82 ( .A(reset), .ZN(n3) );
endmodule


module NRegister_N32_33 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, net108194, net108195, net108196, net108197,
         net108198, net108199, net108200, net108201, net108202, net108203,
         net108204, net108205, net108206, net108207, net108208, net108209,
         net108210, net108211, net108212, net108213, net108214, net108215,
         net108216, net108217, net108218, net108219, net108220, net108221,
         net108222, net108223, net108224, net108225, n35, n36, n37, n38, n39,
         n40, n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53,
         n54, n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67,
         n70, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n44), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n44), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n44), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n46), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n44), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n46), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n46), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n46), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n44), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n46), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n46), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n46), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n46), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n45), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n45), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n45), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n45), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n45), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n45), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n45), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n45), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n45), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n44), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n44), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n44), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n44), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n44), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n44), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n44), .Q(data_out[0]), 
        .QN(net108194) );
  INV_X1 U3 ( .A(n43), .ZN(n36) );
  INV_X1 U4 ( .A(n43), .ZN(n35) );
  BUF_X1 U5 ( .A(n90), .Z(n39) );
  BUF_X1 U6 ( .A(n90), .Z(n40) );
  BUF_X1 U7 ( .A(n90), .Z(n42) );
  BUF_X1 U8 ( .A(n90), .Z(n37) );
  BUF_X1 U9 ( .A(n90), .Z(n38) );
  BUF_X1 U10 ( .A(n90), .Z(n41) );
  BUF_X1 U11 ( .A(n90), .Z(n43) );
  BUF_X1 U12 ( .A(n3), .Z(n45) );
  BUF_X1 U13 ( .A(n3), .Z(n44) );
  BUF_X1 U14 ( .A(n3), .Z(n46) );
  OAI22_X1 U15 ( .A1(n38), .A2(n83), .B1(net108194), .B2(n36), .ZN(n34) );
  INV_X1 U16 ( .A(data_in[0]), .ZN(n83) );
  OAI22_X1 U17 ( .A1(n38), .A2(n82), .B1(net108195), .B2(n35), .ZN(n33) );
  INV_X1 U18 ( .A(data_in[1]), .ZN(n82) );
  OAI22_X1 U19 ( .A1(n37), .A2(n89), .B1(net108219), .B2(n36), .ZN(n9) );
  INV_X1 U20 ( .A(data_in[25]), .ZN(n89) );
  OAI22_X1 U21 ( .A1(n37), .A2(n88), .B1(net108220), .B2(n35), .ZN(n8) );
  INV_X1 U22 ( .A(data_in[26]), .ZN(n88) );
  OAI22_X1 U23 ( .A1(n37), .A2(n87), .B1(net108221), .B2(n36), .ZN(n7) );
  INV_X1 U24 ( .A(data_in[27]), .ZN(n87) );
  OAI22_X1 U25 ( .A1(n37), .A2(n86), .B1(net108222), .B2(n35), .ZN(n6) );
  INV_X1 U26 ( .A(data_in[28]), .ZN(n86) );
  OAI22_X1 U27 ( .A1(n37), .A2(n85), .B1(net108223), .B2(n36), .ZN(n5) );
  INV_X1 U28 ( .A(data_in[29]), .ZN(n85) );
  OAI22_X1 U29 ( .A1(n38), .A2(n84), .B1(net108224), .B2(n35), .ZN(n4) );
  INV_X1 U30 ( .A(data_in[30]), .ZN(n84) );
  OAI22_X1 U31 ( .A1(n38), .A2(n81), .B1(net108196), .B2(n36), .ZN(n32) );
  INV_X1 U32 ( .A(data_in[2]), .ZN(n81) );
  OAI22_X1 U33 ( .A1(n38), .A2(n80), .B1(net108197), .B2(n36), .ZN(n31) );
  INV_X1 U34 ( .A(data_in[3]), .ZN(n80) );
  OAI22_X1 U35 ( .A1(n39), .A2(n70), .B1(net108198), .B2(n36), .ZN(n30) );
  INV_X1 U36 ( .A(data_in[4]), .ZN(n70) );
  OAI22_X1 U37 ( .A1(n39), .A2(n67), .B1(net108199), .B2(n36), .ZN(n29) );
  INV_X1 U38 ( .A(data_in[5]), .ZN(n67) );
  OAI22_X1 U39 ( .A1(n39), .A2(n66), .B1(net108200), .B2(n36), .ZN(n28) );
  INV_X1 U40 ( .A(data_in[6]), .ZN(n66) );
  OAI22_X1 U41 ( .A1(n39), .A2(n65), .B1(net108201), .B2(n36), .ZN(n27) );
  INV_X1 U42 ( .A(data_in[7]), .ZN(n65) );
  OAI22_X1 U43 ( .A1(n39), .A2(n64), .B1(net108202), .B2(n36), .ZN(n26) );
  INV_X1 U44 ( .A(data_in[8]), .ZN(n64) );
  OAI22_X1 U45 ( .A1(n40), .A2(n63), .B1(net108203), .B2(n36), .ZN(n25) );
  INV_X1 U46 ( .A(data_in[9]), .ZN(n63) );
  OAI22_X1 U47 ( .A1(n40), .A2(n62), .B1(net108204), .B2(n36), .ZN(n24) );
  INV_X1 U48 ( .A(data_in[10]), .ZN(n62) );
  OAI22_X1 U49 ( .A1(n40), .A2(n61), .B1(net108205), .B2(n36), .ZN(n23) );
  INV_X1 U50 ( .A(data_in[11]), .ZN(n61) );
  OAI22_X1 U51 ( .A1(n40), .A2(n60), .B1(net108206), .B2(n36), .ZN(n22) );
  INV_X1 U52 ( .A(data_in[12]), .ZN(n60) );
  OAI22_X1 U53 ( .A1(n40), .A2(n59), .B1(net108207), .B2(n36), .ZN(n21) );
  INV_X1 U54 ( .A(data_in[13]), .ZN(n59) );
  OAI22_X1 U55 ( .A1(n41), .A2(n58), .B1(net108208), .B2(n35), .ZN(n20) );
  INV_X1 U56 ( .A(data_in[14]), .ZN(n58) );
  OAI22_X1 U57 ( .A1(n41), .A2(n56), .B1(net108209), .B2(n35), .ZN(n19) );
  INV_X1 U58 ( .A(data_in[15]), .ZN(n56) );
  OAI22_X1 U59 ( .A1(n41), .A2(n55), .B1(net108210), .B2(n35), .ZN(n18) );
  INV_X1 U60 ( .A(data_in[16]), .ZN(n55) );
  OAI22_X1 U61 ( .A1(n41), .A2(n54), .B1(net108211), .B2(n35), .ZN(n17) );
  INV_X1 U62 ( .A(data_in[17]), .ZN(n54) );
  OAI22_X1 U63 ( .A1(n42), .A2(n53), .B1(net108212), .B2(n35), .ZN(n16) );
  INV_X1 U64 ( .A(data_in[18]), .ZN(n53) );
  OAI22_X1 U65 ( .A1(n42), .A2(n52), .B1(net108213), .B2(n35), .ZN(n15) );
  INV_X1 U66 ( .A(data_in[19]), .ZN(n52) );
  OAI22_X1 U67 ( .A1(n42), .A2(n51), .B1(net108214), .B2(n35), .ZN(n14) );
  INV_X1 U68 ( .A(data_in[20]), .ZN(n51) );
  OAI22_X1 U69 ( .A1(n42), .A2(n50), .B1(net108215), .B2(n35), .ZN(n13) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n50) );
  OAI22_X1 U71 ( .A1(n42), .A2(n49), .B1(net108216), .B2(n35), .ZN(n12) );
  INV_X1 U72 ( .A(data_in[22]), .ZN(n49) );
  OAI22_X1 U73 ( .A1(n43), .A2(n48), .B1(net108217), .B2(n35), .ZN(n11) );
  INV_X1 U74 ( .A(data_in[23]), .ZN(n48) );
  OAI22_X1 U75 ( .A1(n43), .A2(n47), .B1(net108218), .B2(n35), .ZN(n10) );
  INV_X1 U76 ( .A(data_in[24]), .ZN(n47) );
  OAI22_X1 U77 ( .A1(n41), .A2(n57), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U78 ( .A(data_in[31]), .ZN(n57) );
  NAND2_X1 U79 ( .A1(load), .A2(enable), .ZN(n90) );
  INV_X1 U80 ( .A(reset), .ZN(n3) );
endmodule


module NRegister_N32_32 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108194, net108195, net108196, net108197, net108198,
         net108199, net108200, net108201, net108202, net108203, net108204,
         net108205, net108206, net108207, net108208, net108209, net108210,
         net108211, net108212, net108213, net108214, net108215, net108216,
         net108217, net108218, net108219, net108220, net108221, net108222,
         net108223, net108224, net108225, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n70, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n46), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n46), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n46), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n44), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n46), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n44), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n44), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n44), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n46), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n44), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n44), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n44), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n44), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n44), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n44), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n44), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n44), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n45), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n45), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n45), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n45), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n45), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n45), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n45), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n45), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n45), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n46), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n46), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n46), .Q(data_out[0]), 
        .QN(net108194) );
  BUF_X1 U3 ( .A(n47), .Z(n45) );
  BUF_X1 U4 ( .A(n47), .Z(n44) );
  BUF_X1 U5 ( .A(n47), .Z(n46) );
  INV_X1 U6 ( .A(reset), .ZN(n47) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n92), .Z(n43) );
  BUF_X1 U10 ( .A(n92), .Z(n39) );
  BUF_X1 U11 ( .A(n92), .Z(n40) );
  BUF_X1 U12 ( .A(n92), .Z(n42) );
  BUF_X1 U13 ( .A(n92), .Z(n37) );
  BUF_X1 U14 ( .A(n92), .Z(n38) );
  BUF_X1 U15 ( .A(n92), .Z(n41) );
  OAI22_X1 U16 ( .A1(n38), .A2(n85), .B1(net108194), .B2(n36), .ZN(n34) );
  INV_X1 U17 ( .A(data_in[0]), .ZN(n85) );
  OAI22_X1 U18 ( .A1(n38), .A2(n84), .B1(net108195), .B2(n35), .ZN(n33) );
  INV_X1 U19 ( .A(data_in[1]), .ZN(n84) );
  OAI22_X1 U20 ( .A1(n37), .A2(n91), .B1(net108219), .B2(n36), .ZN(n9) );
  INV_X1 U21 ( .A(data_in[25]), .ZN(n91) );
  OAI22_X1 U22 ( .A1(n37), .A2(n90), .B1(net108220), .B2(n35), .ZN(n8) );
  INV_X1 U23 ( .A(data_in[26]), .ZN(n90) );
  OAI22_X1 U24 ( .A1(n37), .A2(n89), .B1(net108221), .B2(n36), .ZN(n7) );
  INV_X1 U25 ( .A(data_in[27]), .ZN(n89) );
  OAI22_X1 U26 ( .A1(n37), .A2(n88), .B1(net108222), .B2(n35), .ZN(n6) );
  INV_X1 U27 ( .A(data_in[28]), .ZN(n88) );
  OAI22_X1 U28 ( .A1(n37), .A2(n87), .B1(net108223), .B2(n36), .ZN(n5) );
  INV_X1 U29 ( .A(data_in[29]), .ZN(n87) );
  OAI22_X1 U30 ( .A1(n38), .A2(n86), .B1(net108224), .B2(n35), .ZN(n4) );
  INV_X1 U31 ( .A(data_in[30]), .ZN(n86) );
  OAI22_X1 U32 ( .A1(n38), .A2(n83), .B1(net108196), .B2(n36), .ZN(n32) );
  INV_X1 U33 ( .A(data_in[2]), .ZN(n83) );
  OAI22_X1 U34 ( .A1(n38), .A2(n82), .B1(net108197), .B2(n36), .ZN(n31) );
  INV_X1 U35 ( .A(data_in[3]), .ZN(n82) );
  OAI22_X1 U36 ( .A1(n39), .A2(n81), .B1(net108198), .B2(n36), .ZN(n30) );
  INV_X1 U37 ( .A(data_in[4]), .ZN(n81) );
  OAI22_X1 U38 ( .A1(n39), .A2(n70), .B1(net108199), .B2(n36), .ZN(n29) );
  INV_X1 U39 ( .A(data_in[5]), .ZN(n70) );
  OAI22_X1 U40 ( .A1(n39), .A2(n67), .B1(net108200), .B2(n36), .ZN(n28) );
  INV_X1 U41 ( .A(data_in[6]), .ZN(n67) );
  OAI22_X1 U42 ( .A1(n39), .A2(n66), .B1(net108201), .B2(n36), .ZN(n27) );
  INV_X1 U43 ( .A(data_in[7]), .ZN(n66) );
  OAI22_X1 U44 ( .A1(n39), .A2(n65), .B1(net108202), .B2(n36), .ZN(n26) );
  INV_X1 U45 ( .A(data_in[8]), .ZN(n65) );
  OAI22_X1 U46 ( .A1(n40), .A2(n64), .B1(net108203), .B2(n36), .ZN(n25) );
  INV_X1 U47 ( .A(data_in[9]), .ZN(n64) );
  OAI22_X1 U48 ( .A1(n40), .A2(n63), .B1(net108204), .B2(n36), .ZN(n24) );
  INV_X1 U49 ( .A(data_in[10]), .ZN(n63) );
  OAI22_X1 U50 ( .A1(n40), .A2(n62), .B1(net108205), .B2(n36), .ZN(n23) );
  INV_X1 U51 ( .A(data_in[11]), .ZN(n62) );
  OAI22_X1 U52 ( .A1(n40), .A2(n61), .B1(net108206), .B2(n36), .ZN(n22) );
  INV_X1 U53 ( .A(data_in[12]), .ZN(n61) );
  OAI22_X1 U54 ( .A1(n40), .A2(n60), .B1(net108207), .B2(n36), .ZN(n21) );
  INV_X1 U55 ( .A(data_in[13]), .ZN(n60) );
  OAI22_X1 U56 ( .A1(n41), .A2(n59), .B1(net108208), .B2(n35), .ZN(n20) );
  INV_X1 U57 ( .A(data_in[14]), .ZN(n59) );
  OAI22_X1 U58 ( .A1(n41), .A2(n57), .B1(net108209), .B2(n35), .ZN(n19) );
  INV_X1 U59 ( .A(data_in[15]), .ZN(n57) );
  OAI22_X1 U60 ( .A1(n41), .A2(n56), .B1(net108210), .B2(n35), .ZN(n18) );
  INV_X1 U61 ( .A(data_in[16]), .ZN(n56) );
  OAI22_X1 U62 ( .A1(n41), .A2(n55), .B1(net108211), .B2(n35), .ZN(n17) );
  INV_X1 U63 ( .A(data_in[17]), .ZN(n55) );
  OAI22_X1 U64 ( .A1(n42), .A2(n54), .B1(net108212), .B2(n35), .ZN(n16) );
  INV_X1 U65 ( .A(data_in[18]), .ZN(n54) );
  OAI22_X1 U66 ( .A1(n42), .A2(n53), .B1(net108213), .B2(n35), .ZN(n15) );
  INV_X1 U67 ( .A(data_in[19]), .ZN(n53) );
  OAI22_X1 U68 ( .A1(n42), .A2(n52), .B1(net108214), .B2(n35), .ZN(n14) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n52) );
  OAI22_X1 U70 ( .A1(n42), .A2(n51), .B1(net108215), .B2(n35), .ZN(n13) );
  INV_X1 U71 ( .A(data_in[21]), .ZN(n51) );
  OAI22_X1 U72 ( .A1(n42), .A2(n50), .B1(net108216), .B2(n35), .ZN(n12) );
  INV_X1 U73 ( .A(data_in[22]), .ZN(n50) );
  OAI22_X1 U74 ( .A1(n43), .A2(n49), .B1(net108217), .B2(n35), .ZN(n11) );
  INV_X1 U75 ( .A(data_in[23]), .ZN(n49) );
  OAI22_X1 U76 ( .A1(n43), .A2(n48), .B1(net108218), .B2(n35), .ZN(n10) );
  INV_X1 U77 ( .A(data_in[24]), .ZN(n48) );
  OAI22_X1 U78 ( .A1(n41), .A2(n58), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U79 ( .A(data_in[31]), .ZN(n58) );
  NAND2_X1 U80 ( .A1(load), .A2(enable), .ZN(n92) );
endmodule


module NRegister_N32_31 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108194, net108195, net108196, net108197, net108198,
         net108199, net108200, net108201, net108202, net108203, net108204,
         net108205, net108206, net108207, net108208, net108209, net108210,
         net108211, net108212, net108213, net108214, net108215, net108216,
         net108217, net108218, net108219, net108220, net108221, net108222,
         net108223, net108224, net108225, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n79), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n79), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n79), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n77), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n79), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n77), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n77), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n77), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n77), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n77), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n77), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n77), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n78), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n78), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n78), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n78), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n78), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n78), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n78), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108194) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108194), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108195), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n70), .B1(net108219), .B2(n36), .ZN(n9) );
  OAI22_X1 U20 ( .A1(n37), .A2(n71), .B1(net108220), .B2(n35), .ZN(n8) );
  OAI22_X1 U21 ( .A1(n37), .A2(n72), .B1(net108221), .B2(n36), .ZN(n7) );
  OAI22_X1 U22 ( .A1(n37), .A2(n73), .B1(net108222), .B2(n35), .ZN(n6) );
  OAI22_X1 U23 ( .A1(n37), .A2(n74), .B1(net108223), .B2(n36), .ZN(n5) );
  OAI22_X1 U24 ( .A1(n38), .A2(n75), .B1(net108224), .B2(n35), .ZN(n4) );
  OAI22_X1 U25 ( .A1(n38), .A2(n46), .B1(net108196), .B2(n36), .ZN(n32) );
  OAI22_X1 U26 ( .A1(n38), .A2(n47), .B1(net108197), .B2(n36), .ZN(n31) );
  OAI22_X1 U27 ( .A1(n39), .A2(n48), .B1(net108198), .B2(n36), .ZN(n30) );
  OAI22_X1 U28 ( .A1(n39), .A2(n49), .B1(net108199), .B2(n36), .ZN(n29) );
  OAI22_X1 U29 ( .A1(n39), .A2(n50), .B1(net108200), .B2(n36), .ZN(n28) );
  OAI22_X1 U30 ( .A1(n39), .A2(n51), .B1(net108201), .B2(n36), .ZN(n27) );
  OAI22_X1 U31 ( .A1(n39), .A2(n52), .B1(net108202), .B2(n36), .ZN(n26) );
  OAI22_X1 U32 ( .A1(n40), .A2(n53), .B1(net108203), .B2(n36), .ZN(n25) );
  OAI22_X1 U33 ( .A1(n40), .A2(n54), .B1(net108204), .B2(n36), .ZN(n24) );
  OAI22_X1 U34 ( .A1(n40), .A2(n55), .B1(net108205), .B2(n36), .ZN(n23) );
  OAI22_X1 U35 ( .A1(n40), .A2(n56), .B1(net108206), .B2(n36), .ZN(n22) );
  OAI22_X1 U36 ( .A1(n40), .A2(n57), .B1(net108207), .B2(n36), .ZN(n21) );
  OAI22_X1 U37 ( .A1(n41), .A2(n58), .B1(net108208), .B2(n35), .ZN(n20) );
  OAI22_X1 U38 ( .A1(n41), .A2(n59), .B1(net108209), .B2(n35), .ZN(n19) );
  OAI22_X1 U39 ( .A1(n41), .A2(n60), .B1(net108210), .B2(n35), .ZN(n18) );
  OAI22_X1 U40 ( .A1(n41), .A2(n61), .B1(net108211), .B2(n35), .ZN(n17) );
  OAI22_X1 U41 ( .A1(n42), .A2(n62), .B1(net108212), .B2(n35), .ZN(n16) );
  OAI22_X1 U42 ( .A1(n42), .A2(n63), .B1(net108213), .B2(n35), .ZN(n15) );
  OAI22_X1 U43 ( .A1(n42), .A2(n64), .B1(net108214), .B2(n35), .ZN(n14) );
  OAI22_X1 U44 ( .A1(n42), .A2(n65), .B1(net108215), .B2(n35), .ZN(n13) );
  OAI22_X1 U45 ( .A1(n42), .A2(n66), .B1(net108216), .B2(n35), .ZN(n12) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108217), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n43), .A2(n69), .B1(net108218), .B2(n35), .ZN(n10) );
  OAI22_X1 U48 ( .A1(n41), .A2(n76), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_24 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108194, net108195, net108196, net108197, net108198,
         net108199, net108200, net108201, net108202, net108203, net108204,
         net108205, net108206, net108207, net108208, net108209, net108210,
         net108211, net108212, net108213, net108214, net108215, net108216,
         net108217, net108218, net108219, net108220, net108221, net108222,
         net108223, net108224, net108225, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n79), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n79), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n79), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n77), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n79), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n77), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n77), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n77), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n77), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n77), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n77), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n77), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n78), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n78), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n78), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n78), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n78), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n78), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n78), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108194) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108194), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108195), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n70), .B1(net108219), .B2(n36), .ZN(n9) );
  OAI22_X1 U20 ( .A1(n37), .A2(n71), .B1(net108220), .B2(n35), .ZN(n8) );
  OAI22_X1 U21 ( .A1(n37), .A2(n72), .B1(net108221), .B2(n36), .ZN(n7) );
  OAI22_X1 U22 ( .A1(n37), .A2(n73), .B1(net108222), .B2(n35), .ZN(n6) );
  OAI22_X1 U23 ( .A1(n37), .A2(n74), .B1(net108223), .B2(n36), .ZN(n5) );
  OAI22_X1 U24 ( .A1(n38), .A2(n75), .B1(net108224), .B2(n35), .ZN(n4) );
  OAI22_X1 U25 ( .A1(n38), .A2(n46), .B1(net108196), .B2(n36), .ZN(n32) );
  OAI22_X1 U26 ( .A1(n38), .A2(n47), .B1(net108197), .B2(n36), .ZN(n31) );
  OAI22_X1 U27 ( .A1(n39), .A2(n48), .B1(net108198), .B2(n36), .ZN(n30) );
  OAI22_X1 U28 ( .A1(n39), .A2(n49), .B1(net108199), .B2(n36), .ZN(n29) );
  OAI22_X1 U29 ( .A1(n39), .A2(n50), .B1(net108200), .B2(n36), .ZN(n28) );
  OAI22_X1 U30 ( .A1(n39), .A2(n51), .B1(net108201), .B2(n36), .ZN(n27) );
  OAI22_X1 U31 ( .A1(n39), .A2(n52), .B1(net108202), .B2(n36), .ZN(n26) );
  OAI22_X1 U32 ( .A1(n40), .A2(n53), .B1(net108203), .B2(n36), .ZN(n25) );
  OAI22_X1 U33 ( .A1(n40), .A2(n54), .B1(net108204), .B2(n36), .ZN(n24) );
  OAI22_X1 U34 ( .A1(n40), .A2(n55), .B1(net108205), .B2(n36), .ZN(n23) );
  OAI22_X1 U35 ( .A1(n40), .A2(n56), .B1(net108206), .B2(n36), .ZN(n22) );
  OAI22_X1 U36 ( .A1(n40), .A2(n57), .B1(net108207), .B2(n36), .ZN(n21) );
  OAI22_X1 U37 ( .A1(n41), .A2(n58), .B1(net108208), .B2(n35), .ZN(n20) );
  OAI22_X1 U38 ( .A1(n41), .A2(n59), .B1(net108209), .B2(n35), .ZN(n19) );
  OAI22_X1 U39 ( .A1(n41), .A2(n60), .B1(net108210), .B2(n35), .ZN(n18) );
  OAI22_X1 U40 ( .A1(n41), .A2(n61), .B1(net108211), .B2(n35), .ZN(n17) );
  OAI22_X1 U41 ( .A1(n42), .A2(n62), .B1(net108212), .B2(n35), .ZN(n16) );
  OAI22_X1 U42 ( .A1(n42), .A2(n63), .B1(net108213), .B2(n35), .ZN(n15) );
  OAI22_X1 U43 ( .A1(n42), .A2(n64), .B1(net108214), .B2(n35), .ZN(n14) );
  OAI22_X1 U44 ( .A1(n42), .A2(n65), .B1(net108215), .B2(n35), .ZN(n13) );
  OAI22_X1 U45 ( .A1(n42), .A2(n66), .B1(net108216), .B2(n35), .ZN(n12) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108217), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n43), .A2(n69), .B1(net108218), .B2(n35), .ZN(n10) );
  OAI22_X1 U48 ( .A1(n41), .A2(n76), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_14 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108194, net108195, net108196, net108197, net108198,
         net108199, net108200, net108201, net108202, net108203, net108204,
         net108205, net108206, net108207, net108208, net108209, net108210,
         net108211, net108212, net108213, net108214, net108215, net108216,
         net108217, net108218, net108219, net108220, net108221, net108222,
         net108223, net108224, net108225, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n79), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n79), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n79), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n77), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n79), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n77), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n77), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n77), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n77), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n77), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n77), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n77), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n78), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n78), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n78), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n78), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n78), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n78), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n78), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108194) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108194), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108195), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n70), .B1(net108219), .B2(n36), .ZN(n9) );
  OAI22_X1 U20 ( .A1(n37), .A2(n71), .B1(net108220), .B2(n35), .ZN(n8) );
  OAI22_X1 U21 ( .A1(n37), .A2(n72), .B1(net108221), .B2(n36), .ZN(n7) );
  OAI22_X1 U22 ( .A1(n37), .A2(n73), .B1(net108222), .B2(n35), .ZN(n6) );
  OAI22_X1 U23 ( .A1(n37), .A2(n74), .B1(net108223), .B2(n36), .ZN(n5) );
  OAI22_X1 U24 ( .A1(n38), .A2(n75), .B1(net108224), .B2(n35), .ZN(n4) );
  OAI22_X1 U25 ( .A1(n38), .A2(n46), .B1(net108196), .B2(n36), .ZN(n32) );
  OAI22_X1 U26 ( .A1(n38), .A2(n47), .B1(net108197), .B2(n36), .ZN(n31) );
  OAI22_X1 U27 ( .A1(n39), .A2(n48), .B1(net108198), .B2(n36), .ZN(n30) );
  OAI22_X1 U28 ( .A1(n39), .A2(n49), .B1(net108199), .B2(n36), .ZN(n29) );
  OAI22_X1 U29 ( .A1(n39), .A2(n50), .B1(net108200), .B2(n36), .ZN(n28) );
  OAI22_X1 U30 ( .A1(n39), .A2(n51), .B1(net108201), .B2(n36), .ZN(n27) );
  OAI22_X1 U31 ( .A1(n39), .A2(n52), .B1(net108202), .B2(n36), .ZN(n26) );
  OAI22_X1 U32 ( .A1(n40), .A2(n53), .B1(net108203), .B2(n36), .ZN(n25) );
  OAI22_X1 U33 ( .A1(n40), .A2(n54), .B1(net108204), .B2(n36), .ZN(n24) );
  OAI22_X1 U34 ( .A1(n40), .A2(n55), .B1(net108205), .B2(n36), .ZN(n23) );
  OAI22_X1 U35 ( .A1(n40), .A2(n56), .B1(net108206), .B2(n36), .ZN(n22) );
  OAI22_X1 U36 ( .A1(n40), .A2(n57), .B1(net108207), .B2(n36), .ZN(n21) );
  OAI22_X1 U37 ( .A1(n41), .A2(n58), .B1(net108208), .B2(n35), .ZN(n20) );
  OAI22_X1 U38 ( .A1(n41), .A2(n59), .B1(net108209), .B2(n35), .ZN(n19) );
  OAI22_X1 U39 ( .A1(n41), .A2(n60), .B1(net108210), .B2(n35), .ZN(n18) );
  OAI22_X1 U40 ( .A1(n41), .A2(n61), .B1(net108211), .B2(n35), .ZN(n17) );
  OAI22_X1 U41 ( .A1(n42), .A2(n62), .B1(net108212), .B2(n35), .ZN(n16) );
  OAI22_X1 U42 ( .A1(n42), .A2(n63), .B1(net108213), .B2(n35), .ZN(n15) );
  OAI22_X1 U43 ( .A1(n42), .A2(n64), .B1(net108214), .B2(n35), .ZN(n14) );
  OAI22_X1 U44 ( .A1(n42), .A2(n65), .B1(net108215), .B2(n35), .ZN(n13) );
  OAI22_X1 U45 ( .A1(n42), .A2(n66), .B1(net108216), .B2(n35), .ZN(n12) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108217), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n43), .A2(n69), .B1(net108218), .B2(n35), .ZN(n10) );
  OAI22_X1 U48 ( .A1(n41), .A2(n76), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module NRegister_N32_5 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108194, net108195, net108196, net108197, net108198,
         net108199, net108200, net108201, net108202, net108203, net108204,
         net108205, net108206, net108207, net108208, net108209, net108210,
         net108211, net108212, net108213, net108214, net108215, net108216,
         net108217, net108218, net108219, net108220, net108221, net108222,
         net108223, net108224, net108225, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n79), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n79), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n79), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n77), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n79), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n77), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n77), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n77), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n79), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n77), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n77), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n77), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n77), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n77), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n77), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n77), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n77), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n78), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n78), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n78), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n78), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n78), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n78), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n78), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n78), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n78), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n78), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n78), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n78), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n79), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n79), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n79), .Q(data_out[0]), 
        .QN(net108194) );
  BUF_X1 U3 ( .A(n80), .Z(n78) );
  BUF_X1 U4 ( .A(n80), .Z(n77) );
  BUF_X1 U5 ( .A(n80), .Z(n79) );
  INV_X1 U6 ( .A(reset), .ZN(n80) );
  INV_X1 U7 ( .A(n43), .ZN(n36) );
  INV_X1 U8 ( .A(n43), .ZN(n35) );
  BUF_X1 U9 ( .A(n81), .Z(n39) );
  BUF_X1 U10 ( .A(n81), .Z(n40) );
  BUF_X1 U11 ( .A(n81), .Z(n42) );
  BUF_X1 U12 ( .A(n81), .Z(n37) );
  BUF_X1 U13 ( .A(n81), .Z(n38) );
  BUF_X1 U14 ( .A(n81), .Z(n41) );
  BUF_X1 U15 ( .A(n81), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n81) );
  OAI22_X1 U17 ( .A1(n38), .A2(n44), .B1(net108194), .B2(n36), .ZN(n34) );
  OAI22_X1 U18 ( .A1(n38), .A2(n45), .B1(net108195), .B2(n35), .ZN(n33) );
  OAI22_X1 U19 ( .A1(n37), .A2(n70), .B1(net108219), .B2(n36), .ZN(n9) );
  OAI22_X1 U20 ( .A1(n37), .A2(n71), .B1(net108220), .B2(n35), .ZN(n8) );
  OAI22_X1 U21 ( .A1(n37), .A2(n72), .B1(net108221), .B2(n36), .ZN(n7) );
  OAI22_X1 U22 ( .A1(n37), .A2(n73), .B1(net108222), .B2(n35), .ZN(n6) );
  OAI22_X1 U23 ( .A1(n37), .A2(n74), .B1(net108223), .B2(n36), .ZN(n5) );
  OAI22_X1 U24 ( .A1(n38), .A2(n75), .B1(net108224), .B2(n35), .ZN(n4) );
  OAI22_X1 U25 ( .A1(n38), .A2(n46), .B1(net108196), .B2(n36), .ZN(n32) );
  OAI22_X1 U26 ( .A1(n38), .A2(n47), .B1(net108197), .B2(n36), .ZN(n31) );
  OAI22_X1 U27 ( .A1(n39), .A2(n48), .B1(net108198), .B2(n36), .ZN(n30) );
  OAI22_X1 U28 ( .A1(n39), .A2(n49), .B1(net108199), .B2(n36), .ZN(n29) );
  OAI22_X1 U29 ( .A1(n39), .A2(n50), .B1(net108200), .B2(n36), .ZN(n28) );
  OAI22_X1 U30 ( .A1(n39), .A2(n51), .B1(net108201), .B2(n36), .ZN(n27) );
  OAI22_X1 U31 ( .A1(n39), .A2(n52), .B1(net108202), .B2(n36), .ZN(n26) );
  OAI22_X1 U32 ( .A1(n40), .A2(n53), .B1(net108203), .B2(n36), .ZN(n25) );
  OAI22_X1 U33 ( .A1(n40), .A2(n54), .B1(net108204), .B2(n36), .ZN(n24) );
  OAI22_X1 U34 ( .A1(n40), .A2(n55), .B1(net108205), .B2(n36), .ZN(n23) );
  OAI22_X1 U35 ( .A1(n40), .A2(n56), .B1(net108206), .B2(n36), .ZN(n22) );
  OAI22_X1 U36 ( .A1(n40), .A2(n57), .B1(net108207), .B2(n36), .ZN(n21) );
  OAI22_X1 U37 ( .A1(n41), .A2(n58), .B1(net108208), .B2(n35), .ZN(n20) );
  OAI22_X1 U38 ( .A1(n41), .A2(n59), .B1(net108209), .B2(n35), .ZN(n19) );
  OAI22_X1 U39 ( .A1(n41), .A2(n60), .B1(net108210), .B2(n35), .ZN(n18) );
  OAI22_X1 U40 ( .A1(n41), .A2(n61), .B1(net108211), .B2(n35), .ZN(n17) );
  OAI22_X1 U41 ( .A1(n42), .A2(n62), .B1(net108212), .B2(n35), .ZN(n16) );
  OAI22_X1 U42 ( .A1(n42), .A2(n63), .B1(net108213), .B2(n35), .ZN(n15) );
  OAI22_X1 U43 ( .A1(n42), .A2(n64), .B1(net108214), .B2(n35), .ZN(n14) );
  OAI22_X1 U44 ( .A1(n42), .A2(n65), .B1(net108215), .B2(n35), .ZN(n13) );
  OAI22_X1 U45 ( .A1(n42), .A2(n66), .B1(net108216), .B2(n35), .ZN(n12) );
  OAI22_X1 U46 ( .A1(n43), .A2(n67), .B1(net108217), .B2(n35), .ZN(n11) );
  OAI22_X1 U47 ( .A1(n43), .A2(n69), .B1(net108218), .B2(n35), .ZN(n10) );
  OAI22_X1 U48 ( .A1(n41), .A2(n76), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U49 ( .A(data_in[0]), .ZN(n44) );
  INV_X1 U50 ( .A(data_in[1]), .ZN(n45) );
  INV_X1 U51 ( .A(data_in[2]), .ZN(n46) );
  INV_X1 U52 ( .A(data_in[3]), .ZN(n47) );
  INV_X1 U53 ( .A(data_in[4]), .ZN(n48) );
  INV_X1 U54 ( .A(data_in[5]), .ZN(n49) );
  INV_X1 U55 ( .A(data_in[6]), .ZN(n50) );
  INV_X1 U56 ( .A(data_in[7]), .ZN(n51) );
  INV_X1 U57 ( .A(data_in[8]), .ZN(n52) );
  INV_X1 U58 ( .A(data_in[9]), .ZN(n53) );
  INV_X1 U59 ( .A(data_in[10]), .ZN(n54) );
  INV_X1 U60 ( .A(data_in[11]), .ZN(n55) );
  INV_X1 U61 ( .A(data_in[12]), .ZN(n56) );
  INV_X1 U62 ( .A(data_in[13]), .ZN(n57) );
  INV_X1 U63 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U64 ( .A(data_in[15]), .ZN(n59) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n60) );
  INV_X1 U66 ( .A(data_in[17]), .ZN(n61) );
  INV_X1 U67 ( .A(data_in[18]), .ZN(n62) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n63) );
  INV_X1 U69 ( .A(data_in[20]), .ZN(n64) );
  INV_X1 U70 ( .A(data_in[21]), .ZN(n65) );
  INV_X1 U71 ( .A(data_in[22]), .ZN(n66) );
  INV_X1 U72 ( .A(data_in[23]), .ZN(n67) );
  INV_X1 U73 ( .A(data_in[24]), .ZN(n69) );
  INV_X1 U74 ( .A(data_in[25]), .ZN(n70) );
  INV_X1 U75 ( .A(data_in[26]), .ZN(n71) );
  INV_X1 U76 ( .A(data_in[27]), .ZN(n72) );
  INV_X1 U77 ( .A(data_in[28]), .ZN(n73) );
  INV_X1 U78 ( .A(data_in[29]), .ZN(n74) );
  INV_X1 U79 ( .A(data_in[30]), .ZN(n75) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n76) );
endmodule


module Reg1Bit_22 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n5), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n4), .ZN(n2) );
  INV_X1 U4 ( .A(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U6 ( .A(data_in), .ZN(n4) );
  INV_X1 U7 ( .A(reset), .ZN(n5) );
endmodule


module Reg1Bit_21 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n4), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n5), .ZN(n2) );
  INV_X1 U4 ( .A(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U6 ( .A(data_in), .ZN(n5) );
  INV_X1 U7 ( .A(reset), .ZN(n4) );
endmodule


module Reg1Bit_20 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n4), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n5), .ZN(n2) );
  INV_X1 U4 ( .A(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U6 ( .A(data_in), .ZN(n5) );
  INV_X1 U7 ( .A(reset), .ZN(n4) );
endmodule


module Reg1Bit_19 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n4), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n5), .ZN(n2) );
  INV_X1 U4 ( .A(data_in), .ZN(n5) );
  INV_X1 U5 ( .A(n8), .ZN(n9) );
  NAND2_X1 U6 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U7 ( .A(reset), .ZN(n4) );
endmodule


module Reg1Bit_18 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n4), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n5), .ZN(n2) );
  INV_X1 U4 ( .A(data_in), .ZN(n5) );
  INV_X1 U5 ( .A(n8), .ZN(n9) );
  NAND2_X1 U6 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U7 ( .A(reset), .ZN(n4) );
endmodule


module Reg1Bit_17 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n4), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n5), .ZN(n2) );
  INV_X1 U4 ( .A(data_in), .ZN(n5) );
  INV_X1 U5 ( .A(n8), .ZN(n9) );
  NAND2_X1 U6 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U7 ( .A(reset), .ZN(n4) );
endmodule


module Reg1Bit_16 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, n3, net106835, n4, n5, n7;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n3), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n7), .B1(n5), .B2(n4), .ZN(n2) );
  INV_X1 U4 ( .A(data_in), .ZN(n4) );
  INV_X1 U5 ( .A(n5), .ZN(n7) );
  NAND2_X1 U6 ( .A1(load), .A2(enable), .ZN(n5) );
  INV_X1 U7 ( .A(reset), .ZN(n3) );
endmodule


module Reg1Bit_15 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, n3, net106835, n4, n5, n7;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n3), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n7), .B1(n5), .B2(n4), .ZN(n2) );
  INV_X1 U4 ( .A(data_in), .ZN(n4) );
  INV_X1 U5 ( .A(n5), .ZN(n7) );
  NAND2_X1 U6 ( .A1(load), .A2(enable), .ZN(n5) );
  INV_X1 U7 ( .A(reset), .ZN(n3) );
endmodule


module Reg1Bit_14 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n5), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n4), .ZN(n2) );
  INV_X1 U4 ( .A(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U6 ( .A(data_in), .ZN(n4) );
  INV_X1 U7 ( .A(reset), .ZN(n5) );
endmodule


module Reg1Bit_13 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n5), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n4), .ZN(n2) );
  INV_X1 U4 ( .A(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U6 ( .A(data_in), .ZN(n4) );
  INV_X1 U7 ( .A(reset), .ZN(n5) );
endmodule


module Reg1Bit_12 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n4), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n5), .ZN(n2) );
  INV_X1 U4 ( .A(data_in), .ZN(n5) );
  INV_X1 U5 ( .A(n8), .ZN(n9) );
  NAND2_X1 U6 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U7 ( .A(reset), .ZN(n4) );
endmodule


module Reg1Bit_11 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n4), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n5), .ZN(n2) );
  INV_X1 U4 ( .A(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U6 ( .A(data_in), .ZN(n5) );
  INV_X1 U7 ( .A(reset), .ZN(n4) );
endmodule


module Reg1Bit_10 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n5), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n4), .ZN(n2) );
  INV_X1 U4 ( .A(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U6 ( .A(data_in), .ZN(n4) );
  INV_X1 U7 ( .A(reset), .ZN(n5) );
endmodule


module Reg1Bit_9 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n5), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n4), .ZN(n2) );
  INV_X1 U4 ( .A(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U6 ( .A(data_in), .ZN(n4) );
  INV_X1 U7 ( .A(reset), .ZN(n5) );
endmodule


module Reg1Bit_8 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, n3, net106835, n4, n5, n7;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n3), .Q(data_out), .QN(
        net106835) );
  INV_X1 U3 ( .A(reset), .ZN(n3) );
  OAI22_X1 U4 ( .A1(net106835), .A2(n7), .B1(n5), .B2(n4), .ZN(n2) );
  INV_X1 U5 ( .A(n5), .ZN(n7) );
  NAND2_X1 U6 ( .A1(load), .A2(enable), .ZN(n5) );
  INV_X1 U7 ( .A(data_in), .ZN(n4) );
endmodule


module Reg1Bit_7 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n5), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n4), .ZN(n2) );
  INV_X1 U4 ( .A(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U6 ( .A(data_in), .ZN(n4) );
  INV_X1 U7 ( .A(reset), .ZN(n5) );
endmodule


module Reg1Bit_6 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n4), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n5), .ZN(n2) );
  INV_X1 U4 ( .A(data_in), .ZN(n5) );
  INV_X1 U5 ( .A(n8), .ZN(n9) );
  NAND2_X1 U6 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U7 ( .A(reset), .ZN(n4) );
endmodule


module Reg1Bit_5 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n4), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n5), .ZN(n2) );
  INV_X1 U4 ( .A(data_in), .ZN(n5) );
  INV_X1 U5 ( .A(n8), .ZN(n9) );
  NAND2_X1 U6 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U7 ( .A(reset), .ZN(n4) );
endmodule


module Reg1Bit_4 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n4), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n5), .ZN(n2) );
  INV_X1 U4 ( .A(data_in), .ZN(n5) );
  INV_X1 U5 ( .A(n8), .ZN(n9) );
  NAND2_X1 U6 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U7 ( .A(reset), .ZN(n4) );
endmodule


module Reg1Bit_3 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n4), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n5), .ZN(n2) );
  INV_X1 U4 ( .A(data_in), .ZN(n5) );
  INV_X1 U5 ( .A(n8), .ZN(n9) );
  NAND2_X1 U6 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U7 ( .A(reset), .ZN(n4) );
endmodule


module Reg1Bit_2 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n4), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n5), .ZN(n2) );
  INV_X1 U4 ( .A(data_in), .ZN(n5) );
  INV_X1 U5 ( .A(n8), .ZN(n9) );
  NAND2_X1 U6 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U7 ( .A(reset), .ZN(n4) );
endmodule


module Reg1Bit_1 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n4, n5, n8, n9;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n4), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n9), .B1(n8), .B2(n5), .ZN(n2) );
  INV_X1 U4 ( .A(n8), .ZN(n9) );
  NAND2_X1 U5 ( .A1(load), .A2(enable), .ZN(n8) );
  INV_X1 U6 ( .A(data_in), .ZN(n5) );
  INV_X1 U7 ( .A(reset), .ZN(n4) );
endmodule


module MUX21_0 ( A, B, S, Y );
  input A, B, S;
  output Y;
  wire   n3, n1;

  INV_X1 U1 ( .A(n3), .ZN(Y) );
  AOI22_X1 U2 ( .A1(A), .A2(n1), .B1(S), .B2(B), .ZN(n3) );
  INV_X1 U3 ( .A(S), .ZN(n1) );
endmodule


module FA_0 ( A, B, Ci, S, Co );
  input A, B, Ci;
  output S, Co;
  wire   n2, n3;

  XOR2_X1 U3 ( .A(Ci), .B(n2), .Z(S) );
  XOR2_X1 U4 ( .A(A), .B(B), .Z(n2) );
  INV_X1 U1 ( .A(n3), .ZN(Co) );
  AOI22_X1 U2 ( .A1(B), .A2(A), .B1(n2), .B2(Ci), .ZN(n3) );
endmodule


module MUX21_GENERIC_N4_0 ( A, B, SEL, Y );
  input [3:0] A;
  input [3:0] B;
  output [3:0] Y;
  input SEL;


  MUX21_0 U_0 ( .A(A[0]), .B(B[0]), .S(SEL), .Y(Y[0]) );
  MUX21_31 U_1 ( .A(A[1]), .B(B[1]), .S(SEL), .Y(Y[1]) );
  MUX21_30 U_2 ( .A(A[2]), .B(B[2]), .S(SEL), .Y(Y[2]) );
  MUX21_29 U_3 ( .A(A[3]), .B(B[3]), .S(SEL), .Y(Y[3]) );
endmodule


module RCA_N4_0 ( A, B, Ci, S, Co );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Ci;
  output Co;

  wire   [3:1] CTMP;

  FA_0 FAI_1 ( .A(A[0]), .B(B[0]), .Ci(Ci), .S(S[0]), .Co(CTMP[1]) );
  FA_63 FAI_2 ( .A(A[1]), .B(B[1]), .Ci(CTMP[1]), .S(S[1]), .Co(CTMP[2]) );
  FA_62 FAI_3 ( .A(A[2]), .B(B[2]), .Ci(CTMP[2]), .S(S[2]), .Co(CTMP[3]) );
  FA_61 FAI_4 ( .A(A[3]), .B(B[3]), .Ci(CTMP[3]), .S(S[3]), .Co(Co) );
endmodule


module ORGate_NX1_N32_2 ( A, B, Y );
  input [31:0] A;
  input [31:0] B;
  output Y;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26;

  NAND2_X1 U1 ( .A1(n21), .A2(n22), .ZN(Y) );
  AND3_X1 U2 ( .A1(n13), .A2(n15), .A3(n24), .ZN(n21) );
  NOR3_X1 U3 ( .A1(n1), .A2(n3), .A3(n4), .ZN(n22) );
  AND3_X1 U4 ( .A1(n19), .A2(n20), .A3(n17), .ZN(n23) );
  AND2_X1 U5 ( .A1(n14), .A2(n16), .ZN(n24) );
  OR3_X1 U6 ( .A1(A[28]), .A2(A[29]), .A3(A[30]), .ZN(n25) );
  NOR4_X1 U7 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n15) );
  NAND2_X1 U8 ( .A1(n18), .A2(n23), .ZN(n1) );
  NOR2_X1 U9 ( .A1(A[2]), .A2(n25), .ZN(n18) );
  NOR4_X1 U10 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n16) );
  NOR4_X1 U11 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n14) );
  NOR4_X1 U12 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n19) );
  OR3_X1 U13 ( .A1(A[10]), .A2(A[11]), .A3(A[12]), .ZN(n26) );
  NOR4_X1 U14 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n20) );
  NOR4_X1 U15 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n17) );
  NAND4_X1 U16 ( .A1(n5), .A2(n6), .A3(n7), .A4(n8), .ZN(n4) );
  NAND4_X1 U17 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .ZN(n3) );
  NOR4_X1 U18 ( .A1(B[9]), .A2(B[8]), .A3(B[7]), .A4(B[6]), .ZN(n12) );
  NOR4_X1 U19 ( .A1(B[23]), .A2(B[22]), .A3(B[21]), .A4(B[20]), .ZN(n8) );
  NOR4_X1 U20 ( .A1(B[5]), .A2(B[4]), .A3(B[3]), .A4(B[31]), .ZN(n11) );
  NOR4_X1 U21 ( .A1(B[1]), .A2(B[19]), .A3(B[18]), .A4(B[17]), .ZN(n7) );
  NOR4_X1 U22 ( .A1(B[30]), .A2(B[2]), .A3(B[29]), .A4(B[28]), .ZN(n10) );
  NOR4_X1 U23 ( .A1(B[16]), .A2(B[15]), .A3(B[14]), .A4(B[13]), .ZN(n6) );
  NOR4_X1 U24 ( .A1(B[27]), .A2(B[26]), .A3(B[25]), .A4(B[24]), .ZN(n9) );
  NOR4_X1 U25 ( .A1(B[12]), .A2(B[11]), .A3(B[10]), .A4(B[0]), .ZN(n5) );
  NOR2_X1 U26 ( .A1(A[0]), .A2(n26), .ZN(n13) );
endmodule


module CarrySelectBlock_N4_0 ( A, B, Cin, S );
  input [3:0] A;
  input [3:0] B;
  output [3:0] S;
  input Cin;

  wire   [3:0] sum1;
  wire   [3:0] sum2;

  RCA_N4_0 rca1 ( .A(A), .B(B), .Ci(1'b0), .S(sum1) );
  RCA_N4_15 rca2 ( .A(A), .B(B), .Ci(1'b1), .S(sum2) );
  MUX21_GENERIC_N4_0 mux ( .A(sum1), .B(sum2), .SEL(Cin), .Y(S) );
endmodule


module GeneralPropagate_0 ( G_ik, P_ik, G_km1_j, P_km1_j, G_ij, P_ij );
  input G_ik, P_ik, G_km1_j, P_km1_j;
  output G_ij, P_ij;
  wire   n2;

  AND2_X1 U1 ( .A1(P_km1_j), .A2(P_ik), .ZN(P_ij) );
  INV_X1 U2 ( .A(n2), .ZN(G_ij) );
  AOI21_X1 U3 ( .B1(G_km1_j), .B2(P_ik), .A(G_ik), .ZN(n2) );
endmodule


module Multiplier_NBIT_DATA32_DW01_add_1 ( A, B, CI, SUM, CO );
  input [61:0] A;
  input [61:0] B;
  output [61:0] SUM;
  input CI;
  output CO;
  wire   \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] , \A[23] ,
         \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] , \A[16] ,
         \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] , \A[8] ,
         \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] , \A[0] , n1,
         n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n30, n31, n32, n34,
         n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48,
         n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62,
         n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76,
         n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90,
         n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103,
         n104, n105, n106, n107, n108, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n148, n149,
         n150, n152, n153, n154, n155, n156, n157, n158, n159, n160, n161,
         n162, n163, n164, n165, n166, n167, n168, n169, n171, n172, n173,
         n174, n175, n176, n177, n178, n179, n180, n181, n182, n183, n184,
         n185, n186, n187, n188, n189, n190, n191, n192, n193, n194, n195,
         n196, n197, n198, n199, n200, n201, n202, n203, n204, n205, n206,
         n207, n208, n209, n210;
  assign SUM[29] = \A[29] ;
  assign \A[29]  = A[29];
  assign SUM[28] = \A[28] ;
  assign \A[28]  = A[28];
  assign SUM[27] = \A[27] ;
  assign \A[27]  = A[27];
  assign SUM[26] = \A[26] ;
  assign \A[26]  = A[26];
  assign SUM[25] = \A[25] ;
  assign \A[25]  = A[25];
  assign SUM[24] = \A[24] ;
  assign \A[24]  = A[24];
  assign SUM[23] = \A[23] ;
  assign \A[23]  = A[23];
  assign SUM[22] = \A[22] ;
  assign \A[22]  = A[22];
  assign SUM[21] = \A[21] ;
  assign \A[21]  = A[21];
  assign SUM[20] = \A[20] ;
  assign \A[20]  = A[20];
  assign SUM[19] = \A[19] ;
  assign \A[19]  = A[19];
  assign SUM[18] = \A[18] ;
  assign \A[18]  = A[18];
  assign SUM[17] = \A[17] ;
  assign \A[17]  = A[17];
  assign SUM[16] = \A[16] ;
  assign \A[16]  = A[16];
  assign SUM[15] = \A[15] ;
  assign \A[15]  = A[15];
  assign SUM[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2_X1 U6 ( .A(n207), .B(n7), .Z(SUM[60]) );
  XOR2_X1 U18 ( .A(n185), .B(n17), .Z(SUM[58]) );
  XOR2_X1 U25 ( .A(n202), .B(n23), .Z(SUM[57]) );
  XOR2_X1 U30 ( .A(n186), .B(n27), .Z(SUM[56]) );
  XOR2_X1 U42 ( .A(n37), .B(n200), .Z(SUM[54]) );
  XOR2_X1 U49 ( .A(n201), .B(n43), .Z(SUM[53]) );
  XOR2_X1 U54 ( .A(n47), .B(n198), .Z(SUM[52]) );
  XOR2_X1 U61 ( .A(n204), .B(n53), .Z(SUM[51]) );
  XOR2_X1 U66 ( .A(n178), .B(n57), .Z(SUM[50]) );
  XOR2_X1 U73 ( .A(n192), .B(n63), .Z(SUM[49]) );
  XOR2_X1 U78 ( .A(n180), .B(n67), .Z(SUM[48]) );
  XOR2_X1 U97 ( .A(n92), .B(n94), .Z(SUM[46]) );
  XOR2_X1 U109 ( .A(n98), .B(n100), .Z(SUM[44]) );
  XOR2_X1 U119 ( .A(n115), .B(n116), .Z(SUM[43]) );
  XOR2_X1 U126 ( .A(n117), .B(n119), .Z(SUM[42]) );
  XOR2_X1 U155 ( .A(n139), .B(n140), .Z(SUM[38]) );
  XOR2_X1 U160 ( .A(n142), .B(n141), .Z(SUM[37]) );
  XOR2_X1 U167 ( .A(n1), .B(n146), .Z(SUM[36]) );
  XOR2_X1 U178 ( .A(n161), .B(n162), .Z(SUM[35]) );
  XOR2_X1 U185 ( .A(n163), .B(n165), .Z(SUM[34]) );
  XOR2_X1 U190 ( .A(n167), .B(n166), .Z(SUM[33]) );
  XOR2_X1 U197 ( .A(n193), .B(n171), .Z(SUM[32]) );
  XOR2_X1 U203 ( .A(n205), .B(n175), .Z(SUM[31]) );
  NOR4_X2 U147 ( .A1(n125), .A2(n134), .A3(n131), .A4(n135), .ZN(n84) );
  NOR2_X2 U157 ( .A1(B[38]), .A2(A[38]), .ZN(n134) );
  NOR2_X2 U166 ( .A1(B[37]), .A2(A[37]), .ZN(n131) );
  CLKBUF_X1 U2 ( .A(n197), .Z(n178) );
  NOR2_X1 U3 ( .A1(B[41]), .A2(A[41]), .ZN(n109) );
  NOR2_X1 U4 ( .A1(B[36]), .A2(A[36]), .ZN(n135) );
  NOR2_X1 U5 ( .A1(B[39]), .A2(A[39]), .ZN(n125) );
  NOR2_X1 U7 ( .A1(B[44]), .A2(A[44]), .ZN(n99) );
  AND2_X1 U8 ( .A1(B[44]), .A2(A[44]), .ZN(n80) );
  NOR2_X1 U9 ( .A1(B[51]), .A2(A[51]), .ZN(n51) );
  INV_X1 U10 ( .A(n187), .ZN(n164) );
  BUF_X1 U11 ( .A(n189), .Z(n179) );
  CLKBUF_X1 U12 ( .A(n65), .Z(n180) );
  CLKBUF_X1 U13 ( .A(n85), .Z(n181) );
  XNOR2_X1 U14 ( .A(B[61]), .B(A[61]), .ZN(n182) );
  CLKBUF_X1 U15 ( .A(n159), .Z(n183) );
  XNOR2_X1 U16 ( .A(n203), .B(n184), .ZN(SUM[55]) );
  OR2_X1 U17 ( .A1(n30), .A2(n31), .ZN(n184) );
  AOI21_X1 U19 ( .B1(n202), .B2(n18), .A(n20), .ZN(n185) );
  AND2_X1 U20 ( .A1(n153), .A2(n191), .ZN(n86) );
  AOI21_X1 U21 ( .B1(n194), .B2(n28), .A(n30), .ZN(n186) );
  OR2_X2 U22 ( .A1(B[34]), .A2(A[34]), .ZN(n187) );
  XNOR2_X1 U23 ( .A(n208), .B(n188), .ZN(SUM[59]) );
  OR2_X1 U24 ( .A1(n10), .A2(n11), .ZN(n188) );
  OR2_X1 U26 ( .A1(A[33]), .A2(B[33]), .ZN(n189) );
  OAI21_X1 U27 ( .B1(n197), .B2(n54), .A(n56), .ZN(n190) );
  NOR3_X1 U28 ( .A1(n150), .A2(n196), .A3(n148), .ZN(n191) );
  NOR2_X1 U29 ( .A1(A[32]), .A2(B[32]), .ZN(n148) );
  OAI21_X1 U31 ( .B1(n180), .B2(n64), .A(n66), .ZN(n192) );
  OAI21_X1 U32 ( .B1(n172), .B2(n205), .A(n174), .ZN(n193) );
  OAI21_X1 U33 ( .B1(n65), .B2(n64), .A(n66), .ZN(n59) );
  OAI21_X1 U34 ( .B1(n173), .B2(n172), .A(n174), .ZN(n153) );
  OAI21_X1 U35 ( .B1(n35), .B2(n34), .A(n36), .ZN(n194) );
  CLKBUF_X1 U36 ( .A(n172), .Z(n195) );
  OAI21_X1 U37 ( .B1(n55), .B2(n54), .A(n56), .ZN(n49) );
  INV_X1 U38 ( .A(n189), .ZN(n196) );
  AOI21_X1 U39 ( .B1(n192), .B2(n58), .A(n60), .ZN(n197) );
  AOI21_X1 U40 ( .B1(n190), .B2(n48), .A(n50), .ZN(n198) );
  NOR2_X1 U41 ( .A1(B[33]), .A2(A[33]), .ZN(n149) );
  CLKBUF_X1 U43 ( .A(B[30]), .Z(n199) );
  AOI21_X1 U44 ( .B1(n201), .B2(n38), .A(n40), .ZN(n200) );
  OAI21_X1 U45 ( .B1(n44), .B2(n198), .A(n46), .ZN(n201) );
  AOI21_X1 U46 ( .B1(n39), .B2(n38), .A(n40), .ZN(n35) );
  OAI21_X1 U47 ( .B1(n186), .B2(n24), .A(n26), .ZN(n202) );
  OAI21_X1 U48 ( .B1(n34), .B2(n200), .A(n36), .ZN(n203) );
  CLKBUF_X1 U50 ( .A(n190), .Z(n204) );
  OAI21_X1 U51 ( .B1(n25), .B2(n24), .A(n26), .ZN(n19) );
  NAND2_X1 U52 ( .A1(n199), .A2(A[30]), .ZN(n205) );
  AOI21_X1 U53 ( .B1(n202), .B2(n18), .A(n20), .ZN(n206) );
  AOI21_X1 U55 ( .B1(n9), .B2(n8), .A(n10), .ZN(n207) );
  XNOR2_X1 U56 ( .A(n2), .B(n182), .ZN(SUM[61]) );
  OAI21_X1 U57 ( .B1(n206), .B2(n14), .A(n16), .ZN(n208) );
  CLKBUF_X1 U58 ( .A(A[30]), .Z(n209) );
  NAND4_X1 U59 ( .A1(n112), .A2(n107), .A3(n113), .A4(n114), .ZN(n82) );
  AOI21_X1 U60 ( .B1(n1), .B2(n84), .A(n87), .ZN(n101) );
  OAI21_X1 U62 ( .B1(n101), .B2(n82), .A(n83), .ZN(n98) );
  INV_X1 U63 ( .A(n41), .ZN(n38) );
  INV_X1 U64 ( .A(n51), .ZN(n48) );
  NAND2_X1 U65 ( .A1(n12), .A2(n6), .ZN(n7) );
  INV_X1 U67 ( .A(n4), .ZN(n12) );
  NAND2_X1 U68 ( .A1(n22), .A2(n16), .ZN(n17) );
  INV_X1 U69 ( .A(n14), .ZN(n22) );
  NAND2_X1 U70 ( .A1(n32), .A2(n26), .ZN(n27) );
  INV_X1 U71 ( .A(n24), .ZN(n32) );
  NAND2_X1 U72 ( .A1(n42), .A2(n36), .ZN(n37) );
  INV_X1 U74 ( .A(n34), .ZN(n42) );
  NAND2_X1 U75 ( .A1(n52), .A2(n46), .ZN(n47) );
  INV_X1 U76 ( .A(n44), .ZN(n52) );
  NOR2_X1 U77 ( .A1(n20), .A2(n21), .ZN(n23) );
  NOR2_X1 U79 ( .A1(n40), .A2(n41), .ZN(n43) );
  NOR2_X1 U80 ( .A1(n50), .A2(n51), .ZN(n53) );
  AOI21_X1 U81 ( .B1(n194), .B2(n28), .A(n30), .ZN(n25) );
  INV_X1 U82 ( .A(n31), .ZN(n28) );
  AOI21_X1 U83 ( .B1(n19), .B2(n18), .A(n20), .ZN(n15) );
  INV_X1 U84 ( .A(n21), .ZN(n18) );
  AOI21_X1 U85 ( .B1(n157), .B2(n187), .A(n158), .ZN(n155) );
  OAI21_X1 U86 ( .B1(n159), .B2(n149), .A(n160), .ZN(n157) );
  OAI21_X1 U87 ( .B1(n15), .B2(n14), .A(n16), .ZN(n9) );
  AOI21_X1 U88 ( .B1(n59), .B2(n58), .A(n60), .ZN(n55) );
  INV_X1 U89 ( .A(n61), .ZN(n58) );
  AOI21_X1 U90 ( .B1(n9), .B2(n8), .A(n10), .ZN(n5) );
  INV_X1 U91 ( .A(n11), .ZN(n8) );
  AOI21_X1 U92 ( .B1(n78), .B2(n79), .A(n80), .ZN(n76) );
  OAI21_X1 U93 ( .B1(n81), .B2(n82), .A(n83), .ZN(n78) );
  OAI21_X1 U94 ( .B1(n125), .B2(n126), .A(n127), .ZN(n87) );
  AOI21_X1 U95 ( .B1(n128), .B2(n129), .A(n130), .ZN(n126) );
  OAI21_X1 U96 ( .B1(n131), .B2(n132), .A(n133), .ZN(n128) );
  INV_X1 U98 ( .A(n68), .ZN(n65) );
  OAI21_X1 U99 ( .B1(n70), .B2(n69), .A(n71), .ZN(n68) );
  AOI21_X1 U100 ( .B1(n72), .B2(n73), .A(n74), .ZN(n70) );
  OAI21_X1 U101 ( .B1(n76), .B2(n75), .A(n77), .ZN(n72) );
  INV_X1 U102 ( .A(n118), .ZN(n107) );
  INV_X1 U103 ( .A(n109), .ZN(n113) );
  INV_X1 U104 ( .A(n134), .ZN(n129) );
  INV_X1 U105 ( .A(n99), .ZN(n79) );
  INV_X1 U106 ( .A(n154), .ZN(n152) );
  INV_X1 U107 ( .A(n103), .ZN(n112) );
  INV_X1 U108 ( .A(n102), .ZN(n83) );
  OAI21_X1 U110 ( .B1(n103), .B2(n104), .A(n105), .ZN(n102) );
  AOI21_X1 U111 ( .B1(n106), .B2(n107), .A(n108), .ZN(n104) );
  OAI21_X1 U112 ( .B1(n109), .B2(n110), .A(n111), .ZN(n106) );
  INV_X1 U113 ( .A(n123), .ZN(n114) );
  NAND2_X1 U114 ( .A1(n187), .A2(n152), .ZN(n150) );
  AOI21_X1 U115 ( .B1(n79), .B2(n98), .A(n80), .ZN(n95) );
  OAI21_X1 U116 ( .B1(n123), .B2(n101), .A(n110), .ZN(n121) );
  NAND2_X1 U117 ( .A1(n62), .A2(n56), .ZN(n57) );
  INV_X1 U118 ( .A(n54), .ZN(n62) );
  NAND2_X1 U120 ( .A1(n112), .A2(n105), .ZN(n115) );
  AOI21_X1 U121 ( .B1(n117), .B2(n107), .A(n108), .ZN(n116) );
  NAND2_X1 U122 ( .A1(n88), .A2(n66), .ZN(n67) );
  INV_X1 U123 ( .A(n64), .ZN(n88) );
  NAND2_X1 U124 ( .A1(n145), .A2(n133), .ZN(n142) );
  INV_X1 U125 ( .A(n131), .ZN(n145) );
  NAND2_X1 U127 ( .A1(n179), .A2(n160), .ZN(n167) );
  NOR2_X1 U128 ( .A1(n60), .A2(n61), .ZN(n63) );
  NOR2_X1 U129 ( .A1(n74), .A2(n93), .ZN(n94) );
  NOR2_X1 U130 ( .A1(n108), .A2(n118), .ZN(n119) );
  NOR2_X1 U131 ( .A1(n80), .A2(n99), .ZN(n100) );
  NOR2_X1 U132 ( .A1(n158), .A2(n164), .ZN(n165) );
  NOR2_X1 U133 ( .A1(n169), .A2(n148), .ZN(n171) );
  NOR2_X1 U134 ( .A1(n130), .A2(n134), .ZN(n140) );
  NOR2_X1 U135 ( .A1(n144), .A2(n135), .ZN(n146) );
  AOI21_X1 U136 ( .B1(n143), .B2(n1), .A(n144), .ZN(n141) );
  INV_X1 U137 ( .A(n135), .ZN(n143) );
  AOI21_X1 U138 ( .B1(n168), .B2(n193), .A(n169), .ZN(n166) );
  INV_X1 U139 ( .A(n148), .ZN(n168) );
  OAI21_X1 U140 ( .B1(n131), .B2(n141), .A(n133), .ZN(n139) );
  OAI21_X1 U141 ( .B1(n75), .B2(n95), .A(n77), .ZN(n92) );
  OAI21_X1 U142 ( .B1(n196), .B2(n166), .A(n160), .ZN(n163) );
  NAND2_X1 U143 ( .A1(n152), .A2(n156), .ZN(n161) );
  AOI21_X1 U144 ( .B1(n163), .B2(n187), .A(n158), .ZN(n162) );
  XOR2_X1 U145 ( .A(n101), .B(n210), .Z(SUM[40]) );
  NAND2_X1 U146 ( .A1(n110), .A2(n114), .ZN(n210) );
  XNOR2_X1 U148 ( .A(n122), .B(n121), .ZN(SUM[41]) );
  NAND2_X1 U149 ( .A1(n113), .A2(n111), .ZN(n122) );
  XNOR2_X1 U150 ( .A(n95), .B(n96), .ZN(SUM[45]) );
  NOR2_X1 U151 ( .A1(n97), .A2(n75), .ZN(n96) );
  INV_X1 U152 ( .A(n77), .ZN(n97) );
  XNOR2_X1 U153 ( .A(n136), .B(n137), .ZN(SUM[39]) );
  NOR2_X1 U154 ( .A1(n138), .A2(n125), .ZN(n137) );
  AOI21_X1 U156 ( .B1(n129), .B2(n139), .A(n130), .ZN(n136) );
  INV_X1 U158 ( .A(n127), .ZN(n138) );
  XNOR2_X1 U159 ( .A(n89), .B(n90), .ZN(SUM[47]) );
  NOR2_X1 U161 ( .A1(n91), .A2(n69), .ZN(n90) );
  AOI21_X1 U162 ( .B1(n73), .B2(n92), .A(n74), .ZN(n89) );
  INV_X1 U163 ( .A(n71), .ZN(n91) );
  INV_X1 U164 ( .A(n93), .ZN(n73) );
  INV_X1 U165 ( .A(n183), .ZN(n169) );
  INV_X1 U168 ( .A(n132), .ZN(n144) );
  OAI21_X1 U169 ( .B1(n109), .B2(n120), .A(n111), .ZN(n117) );
  INV_X1 U170 ( .A(n121), .ZN(n120) );
  NOR2_X1 U171 ( .A1(B[42]), .A2(A[42]), .ZN(n118) );
  NOR2_X1 U172 ( .A1(B[31]), .A2(A[31]), .ZN(n172) );
  NOR2_X1 U173 ( .A1(B[43]), .A2(A[43]), .ZN(n103) );
  NOR2_X1 U174 ( .A1(B[40]), .A2(A[40]), .ZN(n123) );
  NOR2_X1 U175 ( .A1(B[35]), .A2(A[35]), .ZN(n154) );
  NAND2_X1 U176 ( .A1(A[33]), .A2(B[33]), .ZN(n160) );
  NAND2_X1 U177 ( .A1(B[37]), .A2(A[37]), .ZN(n133) );
  NAND2_X1 U179 ( .A1(B[41]), .A2(A[41]), .ZN(n111) );
  AND2_X1 U180 ( .A1(B[34]), .A2(A[34]), .ZN(n158) );
  AND2_X1 U181 ( .A1(B[38]), .A2(A[38]), .ZN(n130) );
  AND2_X1 U182 ( .A1(B[42]), .A2(A[42]), .ZN(n108) );
  NAND2_X1 U183 ( .A1(B[40]), .A2(A[40]), .ZN(n110) );
  NAND2_X1 U184 ( .A1(B[31]), .A2(A[31]), .ZN(n174) );
  NAND2_X1 U186 ( .A1(B[43]), .A2(A[43]), .ZN(n105) );
  NAND2_X1 U187 ( .A1(A[32]), .A2(B[32]), .ZN(n159) );
  NAND2_X1 U188 ( .A1(B[36]), .A2(A[36]), .ZN(n132) );
  NAND2_X1 U189 ( .A1(B[39]), .A2(A[39]), .ZN(n127) );
  NAND2_X1 U191 ( .A1(B[35]), .A2(A[35]), .ZN(n156) );
  NOR2_X1 U192 ( .A1(B[45]), .A2(A[45]), .ZN(n75) );
  NAND2_X1 U193 ( .A1(n176), .A2(n174), .ZN(n175) );
  INV_X1 U194 ( .A(n195), .ZN(n176) );
  NOR2_X1 U195 ( .A1(B[53]), .A2(A[53]), .ZN(n41) );
  NOR2_X1 U196 ( .A1(B[49]), .A2(A[49]), .ZN(n61) );
  NOR2_X1 U198 ( .A1(B[59]), .A2(A[59]), .ZN(n11) );
  NOR2_X1 U199 ( .A1(B[55]), .A2(A[55]), .ZN(n31) );
  NOR2_X1 U200 ( .A1(B[57]), .A2(A[57]), .ZN(n21) );
  NOR2_X1 U201 ( .A1(B[46]), .A2(A[46]), .ZN(n93) );
  NOR2_X1 U202 ( .A1(B[47]), .A2(A[47]), .ZN(n69) );
  NOR2_X1 U204 ( .A1(B[48]), .A2(A[48]), .ZN(n64) );
  NOR2_X1 U205 ( .A1(B[56]), .A2(A[56]), .ZN(n24) );
  NOR2_X1 U206 ( .A1(B[58]), .A2(A[58]), .ZN(n14) );
  NOR2_X1 U207 ( .A1(B[54]), .A2(A[54]), .ZN(n34) );
  NOR2_X1 U208 ( .A1(B[50]), .A2(A[50]), .ZN(n54) );
  NOR2_X1 U209 ( .A1(B[52]), .A2(A[52]), .ZN(n44) );
  NOR2_X1 U210 ( .A1(B[60]), .A2(A[60]), .ZN(n4) );
  NAND2_X1 U211 ( .A1(B[45]), .A2(A[45]), .ZN(n77) );
  AND2_X1 U212 ( .A1(B[46]), .A2(A[46]), .ZN(n74) );
  NAND2_X1 U213 ( .A1(B[48]), .A2(A[48]), .ZN(n66) );
  NAND2_X1 U214 ( .A1(B[56]), .A2(A[56]), .ZN(n26) );
  NAND2_X1 U215 ( .A1(B[58]), .A2(A[58]), .ZN(n16) );
  NAND2_X1 U216 ( .A1(B[54]), .A2(A[54]), .ZN(n36) );
  NAND2_X1 U217 ( .A1(B[47]), .A2(A[47]), .ZN(n71) );
  NAND2_X1 U218 ( .A1(B[50]), .A2(A[50]), .ZN(n56) );
  NAND2_X1 U219 ( .A1(B[52]), .A2(A[52]), .ZN(n46) );
  NAND2_X1 U220 ( .A1(B[60]), .A2(A[60]), .ZN(n6) );
  AND2_X1 U221 ( .A1(B[49]), .A2(A[49]), .ZN(n60) );
  AND2_X1 U222 ( .A1(B[59]), .A2(A[59]), .ZN(n10) );
  AND2_X1 U223 ( .A1(B[55]), .A2(A[55]), .ZN(n30) );
  AND2_X1 U224 ( .A1(B[57]), .A2(A[57]), .ZN(n20) );
  AND2_X1 U225 ( .A1(B[51]), .A2(A[51]), .ZN(n50) );
  AND2_X1 U226 ( .A1(B[53]), .A2(A[53]), .ZN(n40) );
  INV_X1 U227 ( .A(n177), .ZN(SUM[30]) );
  OAI21_X1 U228 ( .B1(n209), .B2(n199), .A(n205), .ZN(n177) );
  OR2_X1 U229 ( .A1(n181), .A2(n86), .ZN(n1) );
  AOI21_X1 U230 ( .B1(n49), .B2(n48), .A(n50), .ZN(n45) );
  OAI21_X1 U231 ( .B1(n45), .B2(n44), .A(n46), .ZN(n39) );
  OAI21_X1 U232 ( .B1(n5), .B2(n4), .A(n6), .ZN(n2) );
  NAND2_X1 U233 ( .A1(B[30]), .A2(A[30]), .ZN(n173) );
  AOI221_X1 U234 ( .B1(n85), .B2(n84), .C1(n86), .C2(n84), .A(n87), .ZN(n81)
         );
  OAI21_X1 U235 ( .B1(n155), .B2(n154), .A(n156), .ZN(n85) );
endmodule


module Multiplier_NBIT_DATA32_DW01_add_0 ( A, B, CI, SUM, CO );
  input [61:0] A;
  input [61:0] B;
  output [61:0] SUM;
  input CI;
  output CO;
  wire   \A[30] , \A[29] , \A[28] , \A[27] , \A[26] , \A[25] , \A[24] ,
         \A[23] , \A[22] , \A[21] , \A[20] , \A[19] , \A[18] , \A[17] ,
         \A[16] , \A[15] , \A[14] , \A[13] , \A[12] , \A[11] , \A[10] , \A[9] ,
         \A[8] , \A[7] , \A[6] , \A[5] , \A[4] , \A[3] , \A[2] , \A[1] ,
         \A[0] , n1, n2, n44, n48, n54, n55, n57, n58, n64, n68, n90, n91, n93,
         n95, n96, n97, n99, n101, n102, n116, n117, n118, n120, n121, n122,
         n123, n124, n126, n128, n131, n132, n133, n134, n135, n136, n137,
         n138, n140, n141, n142, n143, n144, n145, n147, n148, n153, n161,
         n162, n163, n165, n166, n167, n168, n170, n171, n172, net168728,
         net169229, net169228, net169284, net169295, net169402, net169570,
         net169587, net169631, net169630, net169762, net169854, net169906, n42,
         n41, n17, n15, net169294, n87, n150, n146, n139, n130, n129, n127,
         n63, n52, n51, n62, n61, n53, n49, n47, n46, n45, n40, n59, n56, n50,
         n22, n21, net169790, net169261, n158, n156, n119, n113, n112, n111,
         n110, n109, n106, n104, net169349, n9, n7, n6, n5, n4, n23, n19, n16,
         n13, n12, n11, n10, n94, n92, n75, n72, n70, net169588, n43, n39, n37,
         n36, n35, n33, n32, n31, n30, n29, n27, n26, n25, n20, n89, n74, n71,
         n69, n67, n66, n65, n60, n98, n84, n83, n82, n81, n80, n79, n78, n77,
         n76, n73, n115, n114, n108, n107, n105, n103, n100, net169788,
         net169230, n88, n86, n85, n164, n160, n159, n157, n155, n154, n149,
         n173, n174, n175, n176, n177, n178, n179, n180, n181, n182, n183,
         n184, n185, n186, n187, n188, n189, n190, n191, n192, n193;
  assign SUM[30] = \A[30] ;
  assign \A[30]  = A[30];
  assign SUM[29] = \A[29] ;
  assign \A[29]  = A[29];
  assign SUM[28] = \A[28] ;
  assign \A[28]  = A[28];
  assign SUM[27] = \A[27] ;
  assign \A[27]  = A[27];
  assign SUM[26] = \A[26] ;
  assign \A[26]  = A[26];
  assign SUM[25] = \A[25] ;
  assign \A[25]  = A[25];
  assign SUM[24] = \A[24] ;
  assign \A[24]  = A[24];
  assign SUM[23] = \A[23] ;
  assign \A[23]  = A[23];
  assign SUM[22] = \A[22] ;
  assign \A[22]  = A[22];
  assign SUM[21] = \A[21] ;
  assign \A[21]  = A[21];
  assign SUM[20] = \A[20] ;
  assign \A[20]  = A[20];
  assign SUM[19] = \A[19] ;
  assign \A[19]  = A[19];
  assign SUM[18] = \A[18] ;
  assign \A[18]  = A[18];
  assign SUM[17] = \A[17] ;
  assign \A[17]  = A[17];
  assign SUM[16] = \A[16] ;
  assign \A[16]  = A[16];
  assign SUM[15] = \A[15] ;
  assign \A[15]  = A[15];
  assign SUM[14] = \A[14] ;
  assign \A[14]  = A[14];
  assign SUM[13] = \A[13] ;
  assign \A[13]  = A[13];
  assign SUM[12] = \A[12] ;
  assign \A[12]  = A[12];
  assign SUM[11] = \A[11] ;
  assign \A[11]  = A[11];
  assign SUM[10] = \A[10] ;
  assign \A[10]  = A[10];
  assign SUM[9] = \A[9] ;
  assign \A[9]  = A[9];
  assign SUM[8] = \A[8] ;
  assign \A[8]  = A[8];
  assign SUM[7] = \A[7] ;
  assign \A[7]  = A[7];
  assign SUM[6] = \A[6] ;
  assign \A[6]  = A[6];
  assign SUM[5] = \A[5] ;
  assign \A[5]  = A[5];
  assign SUM[4] = \A[4] ;
  assign \A[4]  = A[4];
  assign SUM[3] = \A[3] ;
  assign \A[3]  = A[3];
  assign SUM[2] = \A[2] ;
  assign \A[2]  = A[2];
  assign SUM[1] = \A[1] ;
  assign \A[1]  = A[1];
  assign SUM[0] = \A[0] ;
  assign \A[0]  = A[0];

  XOR2_X1 U51 ( .A(n178), .B(n44), .Z(SUM[53]) );
  XOR2_X1 U56 ( .A(net169854), .B(n48), .Z(SUM[52]) );
  XOR2_X1 U63 ( .A(net169295), .B(n54), .Z(SUM[51]) );
  XOR2_X1 U68 ( .A(net169631), .B(n58), .Z(SUM[50]) );
  XOR2_X1 U75 ( .A(net169284), .B(n64), .Z(SUM[49]) );
  XOR2_X1 U80 ( .A(net169402), .B(n68), .Z(SUM[48]) );
  XOR2_X1 U99 ( .A(n93), .B(n95), .Z(SUM[46]) );
  XOR2_X1 U111 ( .A(n99), .B(n101), .Z(SUM[44]) );
  XOR2_X1 U121 ( .A(n116), .B(n117), .Z(SUM[43]) );
  XOR2_X1 U128 ( .A(n118), .B(n120), .Z(SUM[42]) );
  XOR2_X1 U157 ( .A(n140), .B(n141), .Z(SUM[38]) );
  XOR2_X1 U162 ( .A(n143), .B(n142), .Z(SUM[37]) );
  XOR2_X1 U169 ( .A(n1), .B(n147), .Z(SUM[36]) );
  XOR2_X1 U179 ( .A(n161), .B(n162), .Z(SUM[35]) );
  XOR2_X1 U186 ( .A(n163), .B(n165), .Z(SUM[34]) );
  XOR2_X1 U191 ( .A(n167), .B(n166), .Z(SUM[33]) );
  XOR2_X1 U198 ( .A(n153), .B(n171), .Z(SUM[32]) );
  XNOR2_X1 U2 ( .A(n181), .B(n173), .ZN(SUM[54]) );
  AND2_X1 U3 ( .A1(n43), .A2(n37), .ZN(n173) );
  XNOR2_X1 U4 ( .A(net169906), .B(n174), .ZN(SUM[55]) );
  OR2_X1 U5 ( .A1(n31), .A2(n32), .ZN(n174) );
  XNOR2_X1 U6 ( .A(n180), .B(n175), .ZN(SUM[56]) );
  AND2_X1 U7 ( .A1(n33), .A2(n27), .ZN(n175) );
  CLKBUF_X1 U8 ( .A(n56), .Z(n177) );
  OAI21_X1 U9 ( .B1(net169587), .B2(n25), .A(n27), .ZN(n176) );
  BUF_X1 U10 ( .A(n176), .Z(n179) );
  INV_X1 U11 ( .A(net169790), .ZN(n154) );
  CLKBUF_X1 U12 ( .A(n189), .Z(n178) );
  CLKBUF_X1 U13 ( .A(net169587), .Z(n180) );
  CLKBUF_X1 U14 ( .A(n192), .Z(n181) );
  OAI21_X1 U15 ( .B1(n177), .B2(n55), .A(n57), .ZN(n182) );
  OAI21_X1 U16 ( .B1(n56), .B2(n55), .A(n57), .ZN(n50) );
  AOI21_X1 U17 ( .B1(n182), .B2(n49), .A(n51), .ZN(n183) );
  XNOR2_X1 U18 ( .A(n179), .B(n184), .ZN(SUM[57]) );
  OR2_X1 U19 ( .A1(n21), .A2(n22), .ZN(n184) );
  XNOR2_X1 U20 ( .A(n191), .B(n185), .ZN(SUM[59]) );
  OR2_X1 U21 ( .A1(n11), .A2(n12), .ZN(n185) );
  XNOR2_X1 U22 ( .A(net169229), .B(n186), .ZN(SUM[58]) );
  AND2_X1 U23 ( .A1(n23), .A2(n17), .ZN(n186) );
  OR2_X1 U24 ( .A1(B[34]), .A2(A[34]), .ZN(n187) );
  CLKBUF_X1 U25 ( .A(n87), .Z(n188) );
  OR2_X1 U26 ( .A1(B[34]), .A2(A[34]), .ZN(net169261) );
  CLKBUF_X1 U27 ( .A(n160), .Z(net169762) );
  OAI21_X1 U28 ( .B1(n183), .B2(n45), .A(n47), .ZN(n189) );
  XNOR2_X1 U29 ( .A(net169630), .B(n190), .ZN(SUM[60]) );
  AND2_X1 U30 ( .A1(n13), .A2(n7), .ZN(n190) );
  OAI21_X1 U31 ( .B1(n46), .B2(n45), .A(n47), .ZN(n40) );
  OAI21_X1 U32 ( .B1(n15), .B2(n16), .A(n17), .ZN(n191) );
  INV_X1 U33 ( .A(B[61]), .ZN(net169349) );
  AOI21_X1 U34 ( .B1(n189), .B2(n39), .A(n41), .ZN(n192) );
  AND2_X1 U35 ( .A1(n86), .A2(n85), .ZN(net169230) );
  NOR3_X1 U36 ( .A1(net169230), .A2(n193), .A3(n88), .ZN(n82) );
  OAI21_X1 U37 ( .B1(n155), .B2(n154), .A(n156), .ZN(n86) );
  CLKBUF_X1 U38 ( .A(n86), .Z(net169294) );
  AOI21_X1 U39 ( .B1(n157), .B2(n187), .A(n158), .ZN(n155) );
  OAI21_X1 U40 ( .B1(n159), .B2(n149), .A(n160), .ZN(n157) );
  NOR2_X1 U41 ( .A1(A[33]), .A2(B[33]), .ZN(n149) );
  NAND2_X1 U42 ( .A1(A[32]), .A2(B[32]), .ZN(n159) );
  NOR4_X1 U43 ( .A1(n126), .A2(n135), .A3(n132), .A4(n136), .ZN(n85) );
  AOI21_X1 U44 ( .B1(n1), .B2(n85), .A(n88), .ZN(n102) );
  AND2_X1 U45 ( .A1(n85), .A2(n87), .ZN(n193) );
  NAND2_X1 U46 ( .A1(net169790), .A2(n156), .ZN(n161) );
  NAND2_X1 U47 ( .A1(net169261), .A2(net169790), .ZN(n150) );
  INV_X1 U48 ( .A(n187), .ZN(n164) );
  AOI21_X1 U49 ( .B1(n163), .B2(n187), .A(n158), .ZN(n162) );
  NOR2_X1 U50 ( .A1(n158), .A2(n164), .ZN(n165) );
  NAND2_X1 U52 ( .A1(A[33]), .A2(B[33]), .ZN(n160) );
  NOR2_X1 U53 ( .A1(B[33]), .A2(A[33]), .ZN(net169570) );
  CLKBUF_X1 U54 ( .A(A[32]), .Z(net169788) );
  NOR2_X1 U55 ( .A1(B[32]), .A2(A[32]), .ZN(n148) );
  AND2_X1 U57 ( .A1(net169788), .A2(B[32]), .ZN(net169228) );
  NOR2_X1 U58 ( .A1(n139), .A2(n126), .ZN(n138) );
  OAI21_X1 U59 ( .B1(n126), .B2(n127), .A(n128), .ZN(n88) );
  NOR2_X1 U60 ( .A1(n131), .A2(n135), .ZN(n141) );
  INV_X1 U61 ( .A(n135), .ZN(n130) );
  OAI21_X1 U62 ( .B1(n132), .B2(n142), .A(n134), .ZN(n140) );
  INV_X1 U64 ( .A(n132), .ZN(n146) );
  OAI21_X1 U65 ( .B1(n132), .B2(n133), .A(n134), .ZN(n129) );
  OAI21_X1 U66 ( .B1(n77), .B2(n76), .A(n78), .ZN(n73) );
  AOI21_X1 U67 ( .B1(n73), .B2(n74), .A(n75), .ZN(n71) );
  AOI21_X1 U69 ( .B1(n79), .B2(n80), .A(n81), .ZN(n77) );
  INV_X1 U70 ( .A(n100), .ZN(n80) );
  AOI21_X1 U71 ( .B1(n80), .B2(n99), .A(n81), .ZN(n96) );
  OAI21_X1 U72 ( .B1(n82), .B2(n83), .A(n84), .ZN(n79) );
  INV_X1 U73 ( .A(n103), .ZN(n84) );
  OAI21_X1 U74 ( .B1(n102), .B2(n83), .A(n84), .ZN(n99) );
  OAI21_X1 U76 ( .B1(n104), .B2(n105), .A(n106), .ZN(n103) );
  AOI21_X1 U77 ( .B1(n107), .B2(n108), .A(n109), .ZN(n105) );
  INV_X1 U78 ( .A(n119), .ZN(n108) );
  NAND4_X1 U79 ( .A1(n113), .A2(n108), .A3(n114), .A4(n115), .ZN(n83) );
  AOI21_X1 U81 ( .B1(n118), .B2(n108), .A(n109), .ZN(n117) );
  OAI21_X1 U82 ( .B1(n110), .B2(n111), .A(n112), .ZN(n107) );
  NOR2_X1 U83 ( .A1(B[45]), .A2(A[45]), .ZN(n76) );
  OAI21_X1 U84 ( .B1(n76), .B2(n96), .A(n78), .ZN(n93) );
  NOR2_X1 U85 ( .A1(n98), .A2(n76), .ZN(n97) );
  NAND2_X1 U86 ( .A1(B[45]), .A2(A[45]), .ZN(n78) );
  INV_X1 U87 ( .A(n78), .ZN(n98) );
  AND2_X1 U88 ( .A1(B[44]), .A2(A[44]), .ZN(n81) );
  NOR2_X1 U89 ( .A1(n81), .A2(n100), .ZN(n101) );
  NOR2_X1 U90 ( .A1(B[44]), .A2(A[44]), .ZN(n100) );
  INV_X1 U91 ( .A(n124), .ZN(n115) );
  NAND2_X1 U92 ( .A1(n111), .A2(n115), .ZN(net168728) );
  INV_X1 U93 ( .A(n110), .ZN(n114) );
  NAND2_X1 U94 ( .A1(n114), .A2(n112), .ZN(n123) );
  INV_X1 U95 ( .A(n104), .ZN(n113) );
  OAI21_X1 U96 ( .B1(n66), .B2(n65), .A(n67), .ZN(n60) );
  AOI21_X1 U97 ( .B1(n60), .B2(n59), .A(n61), .ZN(n56) );
  INV_X1 U98 ( .A(n69), .ZN(n66) );
  CLKBUF_X1 U100 ( .A(n66), .Z(net169402) );
  OAI21_X1 U101 ( .B1(n71), .B2(n70), .A(n72), .ZN(n69) );
  INV_X1 U102 ( .A(n94), .ZN(n74) );
  AOI21_X1 U103 ( .B1(n74), .B2(n93), .A(n75), .ZN(n90) );
  NOR2_X1 U104 ( .A1(B[48]), .A2(A[48]), .ZN(n65) );
  OAI21_X1 U105 ( .B1(n65), .B2(net169402), .A(n67), .ZN(net169284) );
  INV_X1 U106 ( .A(n65), .ZN(n89) );
  NAND2_X1 U107 ( .A1(B[48]), .A2(A[48]), .ZN(n67) );
  NAND2_X1 U108 ( .A1(n89), .A2(n67), .ZN(n68) );
  NOR2_X1 U109 ( .A1(B[47]), .A2(A[47]), .ZN(n70) );
  OAI21_X1 U110 ( .B1(n26), .B2(n25), .A(n27), .ZN(n20) );
  AOI21_X1 U112 ( .B1(n20), .B2(n19), .A(n21), .ZN(n16) );
  AOI21_X1 U113 ( .B1(n30), .B2(n29), .A(n31), .ZN(n26) );
  INV_X1 U114 ( .A(n32), .ZN(n29) );
  AOI21_X1 U115 ( .B1(net169588), .B2(n29), .A(n31), .ZN(net169587) );
  OAI21_X1 U116 ( .B1(n36), .B2(n35), .A(n37), .ZN(n30) );
  NOR2_X1 U117 ( .A1(B[56]), .A2(A[56]), .ZN(n25) );
  INV_X1 U118 ( .A(n25), .ZN(n33) );
  NAND2_X1 U119 ( .A1(B[56]), .A2(A[56]), .ZN(n27) );
  AND2_X1 U120 ( .A1(B[55]), .A2(A[55]), .ZN(n31) );
  NOR2_X1 U122 ( .A1(B[55]), .A2(A[55]), .ZN(n32) );
  AOI21_X1 U123 ( .B1(n40), .B2(n39), .A(n41), .ZN(n36) );
  OAI21_X1 U124 ( .B1(n181), .B2(n35), .A(n37), .ZN(net169906) );
  OAI21_X1 U125 ( .B1(n192), .B2(n35), .A(n37), .ZN(net169588) );
  INV_X1 U126 ( .A(n42), .ZN(n39) );
  NOR2_X1 U127 ( .A1(B[54]), .A2(A[54]), .ZN(n35) );
  INV_X1 U129 ( .A(n35), .ZN(n43) );
  NAND2_X1 U130 ( .A1(B[54]), .A2(A[54]), .ZN(n37) );
  NOR2_X1 U131 ( .A1(n41), .A2(n42), .ZN(n44) );
  NOR2_X1 U132 ( .A1(n92), .A2(n70), .ZN(n91) );
  NAND2_X1 U133 ( .A1(B[47]), .A2(A[47]), .ZN(n72) );
  INV_X1 U134 ( .A(n72), .ZN(n92) );
  AND2_X1 U135 ( .A1(B[46]), .A2(A[46]), .ZN(n75) );
  NOR2_X1 U136 ( .A1(n75), .A2(n94), .ZN(n95) );
  NOR2_X1 U137 ( .A1(B[46]), .A2(A[46]), .ZN(n94) );
  XNOR2_X1 U138 ( .A(n4), .B(net169349), .ZN(SUM[61]) );
  OAI21_X1 U139 ( .B1(n6), .B2(n5), .A(n7), .ZN(n4) );
  AOI21_X1 U140 ( .B1(n10), .B2(n9), .A(n11), .ZN(n6) );
  INV_X1 U141 ( .A(n12), .ZN(n9) );
  AOI21_X1 U142 ( .B1(n191), .B2(n9), .A(n11), .ZN(net169630) );
  NOR2_X1 U143 ( .A1(B[60]), .A2(A[60]), .ZN(n5) );
  INV_X1 U144 ( .A(n5), .ZN(n13) );
  NAND2_X1 U145 ( .A1(B[60]), .A2(A[60]), .ZN(n7) );
  OAI21_X1 U146 ( .B1(n16), .B2(n15), .A(n17), .ZN(n10) );
  INV_X1 U147 ( .A(n22), .ZN(n19) );
  AOI21_X1 U148 ( .B1(n176), .B2(n19), .A(n21), .ZN(net169229) );
  AND2_X1 U149 ( .A1(B[59]), .A2(A[59]), .ZN(n11) );
  NOR2_X1 U150 ( .A1(B[59]), .A2(A[59]), .ZN(n12) );
  INV_X1 U151 ( .A(n15), .ZN(n23) );
  NAND2_X1 U152 ( .A1(n113), .A2(n106), .ZN(n116) );
  NOR2_X1 U153 ( .A1(B[43]), .A2(A[43]), .ZN(n104) );
  NAND2_X1 U154 ( .A1(B[43]), .A2(A[43]), .ZN(n106) );
  AND2_X1 U155 ( .A1(B[42]), .A2(A[42]), .ZN(n109) );
  NOR2_X1 U156 ( .A1(n109), .A2(n119), .ZN(n120) );
  NOR2_X1 U158 ( .A1(B[42]), .A2(A[42]), .ZN(n119) );
  NOR2_X1 U159 ( .A1(B[41]), .A2(A[41]), .ZN(n110) );
  OAI21_X1 U160 ( .B1(n110), .B2(n121), .A(n112), .ZN(n118) );
  NAND2_X1 U161 ( .A1(B[40]), .A2(A[40]), .ZN(n111) );
  OAI21_X1 U163 ( .B1(n124), .B2(n102), .A(n111), .ZN(n122) );
  NAND2_X1 U164 ( .A1(B[41]), .A2(A[41]), .ZN(n112) );
  NAND2_X1 U165 ( .A1(B[35]), .A2(A[35]), .ZN(n156) );
  OR2_X2 U166 ( .A1(B[35]), .A2(A[35]), .ZN(net169790) );
  AND2_X1 U167 ( .A1(B[34]), .A2(A[34]), .ZN(n158) );
  AND2_X1 U168 ( .A1(B[57]), .A2(A[57]), .ZN(n21) );
  NOR2_X1 U170 ( .A1(B[57]), .A2(A[57]), .ZN(n22) );
  CLKBUF_X1 U171 ( .A(n182), .Z(net169295) );
  AOI21_X1 U172 ( .B1(n50), .B2(n49), .A(n51), .ZN(n46) );
  CLKBUF_X1 U173 ( .A(n177), .Z(net169631) );
  INV_X1 U174 ( .A(n62), .ZN(n59) );
  NOR2_X1 U175 ( .A1(B[50]), .A2(A[50]), .ZN(n55) );
  CLKBUF_X1 U176 ( .A(n183), .Z(net169854) );
  INV_X1 U177 ( .A(n52), .ZN(n49) );
  NOR2_X1 U178 ( .A1(B[52]), .A2(A[52]), .ZN(n45) );
  INV_X1 U180 ( .A(n45), .ZN(n53) );
  NAND2_X1 U181 ( .A1(B[52]), .A2(A[52]), .ZN(n47) );
  NAND2_X1 U182 ( .A1(n53), .A2(n47), .ZN(n48) );
  NOR2_X1 U183 ( .A1(n51), .A2(n52), .ZN(n54) );
  AND2_X1 U184 ( .A1(B[49]), .A2(A[49]), .ZN(n61) );
  NOR2_X1 U185 ( .A1(n61), .A2(n62), .ZN(n64) );
  NOR2_X1 U187 ( .A1(B[49]), .A2(A[49]), .ZN(n62) );
  AND2_X1 U188 ( .A1(B[51]), .A2(A[51]), .ZN(n51) );
  NOR2_X1 U189 ( .A1(B[51]), .A2(A[51]), .ZN(n52) );
  INV_X1 U190 ( .A(n55), .ZN(n63) );
  NAND2_X1 U192 ( .A1(n63), .A2(n57), .ZN(n58) );
  AOI21_X1 U193 ( .B1(n129), .B2(n130), .A(n131), .ZN(n127) );
  AOI21_X1 U194 ( .B1(n130), .B2(n140), .A(n131), .ZN(n137) );
  NOR4_X1 U195 ( .A1(n172), .A2(n148), .A3(net169570), .A4(n150), .ZN(n87) );
  OR2_X1 U196 ( .A1(net169294), .A2(n188), .ZN(n1) );
  INV_X1 U197 ( .A(n128), .ZN(n139) );
  INV_X1 U199 ( .A(n133), .ZN(n145) );
  NAND2_X1 U200 ( .A1(n146), .A2(n134), .ZN(n143) );
  NOR2_X1 U201 ( .A1(n145), .A2(n136), .ZN(n147) );
  INV_X1 U202 ( .A(n136), .ZN(n144) );
  NOR2_X1 U203 ( .A1(B[58]), .A2(A[58]), .ZN(n15) );
  NAND2_X1 U204 ( .A1(B[58]), .A2(A[58]), .ZN(n17) );
  AND2_X1 U205 ( .A1(B[53]), .A2(A[53]), .ZN(n41) );
  NOR2_X1 U206 ( .A1(B[53]), .A2(A[53]), .ZN(n42) );
  NAND2_X1 U207 ( .A1(net169762), .A2(n170), .ZN(n167) );
  NOR2_X1 U208 ( .A1(net169228), .A2(n148), .ZN(n171) );
  AOI21_X1 U209 ( .B1(n144), .B2(n1), .A(n145), .ZN(n142) );
  AOI21_X1 U210 ( .B1(n168), .B2(n153), .A(net169228), .ZN(n166) );
  INV_X1 U211 ( .A(n148), .ZN(n168) );
  XOR2_X1 U212 ( .A(n102), .B(net168728), .Z(SUM[40]) );
  XNOR2_X1 U213 ( .A(n123), .B(n122), .ZN(SUM[41]) );
  XNOR2_X1 U214 ( .A(n96), .B(n97), .ZN(SUM[45]) );
  XNOR2_X1 U215 ( .A(n137), .B(n138), .ZN(SUM[39]) );
  XNOR2_X1 U216 ( .A(n90), .B(n91), .ZN(SUM[47]) );
  INV_X1 U217 ( .A(n172), .ZN(n153) );
  INV_X1 U218 ( .A(n122), .ZN(n121) );
  NOR2_X1 U219 ( .A1(B[37]), .A2(A[37]), .ZN(n132) );
  NOR2_X1 U220 ( .A1(B[36]), .A2(A[36]), .ZN(n136) );
  NOR2_X1 U221 ( .A1(B[38]), .A2(A[38]), .ZN(n135) );
  NOR2_X1 U222 ( .A1(B[39]), .A2(A[39]), .ZN(n126) );
  NOR2_X1 U223 ( .A1(B[40]), .A2(A[40]), .ZN(n124) );
  NAND2_X1 U224 ( .A1(B[37]), .A2(A[37]), .ZN(n134) );
  AND2_X1 U225 ( .A1(B[38]), .A2(A[38]), .ZN(n131) );
  NAND2_X1 U226 ( .A1(B[31]), .A2(A[31]), .ZN(n172) );
  NAND2_X1 U227 ( .A1(B[36]), .A2(A[36]), .ZN(n133) );
  NAND2_X1 U228 ( .A1(B[39]), .A2(A[39]), .ZN(n128) );
  NAND2_X1 U229 ( .A1(B[50]), .A2(A[50]), .ZN(n57) );
  AND2_X1 U230 ( .A1(n2), .A2(n172), .ZN(SUM[31]) );
  OR2_X1 U231 ( .A1(B[31]), .A2(A[31]), .ZN(n2) );
  INV_X1 U232 ( .A(net169570), .ZN(n170) );
  OAI21_X1 U233 ( .B1(net169570), .B2(n166), .A(net169762), .ZN(n163) );
endmodule


module XNORGate_NX1_N32 ( A, B, Y );
  input [31:0] A;
  input [31:0] B;
  output Y;
  wire   n1, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n52, n54, n55, n56, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66;

  XOR2_X1 U34 ( .A(n5), .B(n6), .Z(n4) );
  XOR2_X1 U35 ( .A(n7), .B(n8), .Z(n6) );
  XOR2_X1 U36 ( .A(n9), .B(n10), .Z(n8) );
  XOR2_X1 U37 ( .A(n11), .B(n12), .Z(n7) );
  XOR2_X1 U38 ( .A(n13), .B(n14), .Z(n5) );
  XOR2_X1 U39 ( .A(n15), .B(n16), .Z(n14) );
  XOR2_X1 U40 ( .A(n17), .B(n18), .Z(n13) );
  XOR2_X1 U41 ( .A(n19), .B(n20), .Z(n3) );
  XOR2_X1 U42 ( .A(n21), .B(n22), .Z(n20) );
  XOR2_X1 U43 ( .A(n23), .B(n24), .Z(n22) );
  XOR2_X1 U44 ( .A(n25), .B(n26), .Z(n21) );
  XOR2_X1 U45 ( .A(n27), .B(n28), .Z(n19) );
  XOR2_X1 U46 ( .A(n29), .B(n30), .Z(n28) );
  XOR2_X1 U47 ( .A(n31), .B(n32), .Z(n27) );
  XOR2_X1 U49 ( .A(n35), .B(n36), .Z(n34) );
  XOR2_X1 U50 ( .A(n37), .B(n38), .Z(n36) );
  XOR2_X1 U51 ( .A(n39), .B(n40), .Z(n38) );
  XOR2_X1 U52 ( .A(n41), .B(n42), .Z(n37) );
  XOR2_X1 U53 ( .A(n43), .B(n44), .Z(n35) );
  XOR2_X1 U54 ( .A(n45), .B(n46), .Z(n44) );
  XOR2_X1 U55 ( .A(n47), .B(n48), .Z(n43) );
  XOR2_X1 U60 ( .A(n57), .B(n58), .Z(n49) );
  XOR2_X1 U61 ( .A(n59), .B(n60), .Z(n58) );
  XOR2_X1 U62 ( .A(n61), .B(n62), .Z(n57) );
  XOR2_X1 U63 ( .A(A[19]), .B(A[18]), .Z(n62) );
  XNOR2_X1 U1 ( .A(n1), .B(n63), .ZN(Y) );
  XNOR2_X1 U2 ( .A(n3), .B(n4), .ZN(n63) );
  XNOR2_X1 U3 ( .A(A[5]), .B(A[4]), .ZN(n16) );
  XNOR2_X1 U4 ( .A(A[7]), .B(A[6]), .ZN(n15) );
  XNOR2_X1 U5 ( .A(A[27]), .B(A[26]), .ZN(n56) );
  XNOR2_X1 U6 ( .A(A[23]), .B(A[22]), .ZN(n60) );
  XNOR2_X1 U7 ( .A(A[21]), .B(A[20]), .ZN(n46) );
  XNOR2_X1 U8 ( .A(A[15]), .B(A[14]), .ZN(n39) );
  XNOR2_X1 U9 ( .A(A[13]), .B(A[12]), .ZN(n40) );
  XNOR2_X1 U10 ( .A(A[31]), .B(A[30]), .ZN(n9) );
  XNOR2_X1 U11 ( .A(A[29]), .B(A[28]), .ZN(n10) );
  XNOR2_X1 U12 ( .A(A[17]), .B(A[16]), .ZN(n61) );
  XNOR2_X1 U13 ( .A(B[17]), .B(B[16]), .ZN(n55) );
  XNOR2_X1 U14 ( .A(B[31]), .B(B[30]), .ZN(n47) );
  XNOR2_X1 U15 ( .A(B[1]), .B(B[0]), .ZN(n41) );
  XNOR2_X1 U16 ( .A(A[3]), .B(A[2]), .ZN(n42) );
  XNOR2_X1 U17 ( .A(B[11]), .B(B[10]), .ZN(n23) );
  XNOR2_X1 U18 ( .A(A[9]), .B(A[8]), .ZN(n24) );
  XNOR2_X1 U19 ( .A(B[13]), .B(B[12]), .ZN(n29) );
  XNOR2_X1 U20 ( .A(A[11]), .B(A[10]), .ZN(n30) );
  XNOR2_X1 U21 ( .A(B[7]), .B(B[6]), .ZN(n11) );
  XNOR2_X1 U22 ( .A(B[29]), .B(B[28]), .ZN(n12) );
  XNOR2_X1 U23 ( .A(B[9]), .B(B[8]), .ZN(n25) );
  XNOR2_X1 U24 ( .A(B[25]), .B(B[24]), .ZN(n26) );
  XNOR2_X1 U25 ( .A(B[23]), .B(B[22]), .ZN(n48) );
  XNOR2_X1 U26 ( .A(B[27]), .B(B[26]), .ZN(n18) );
  XNOR2_X1 U27 ( .A(B[15]), .B(B[14]), .ZN(n32) );
  XNOR2_X1 U28 ( .A(B[19]), .B(B[18]), .ZN(n59) );
  XNOR2_X1 U29 ( .A(B[21]), .B(B[20]), .ZN(n45) );
  XNOR2_X1 U30 ( .A(B[5]), .B(B[4]), .ZN(n17) );
  XNOR2_X1 U31 ( .A(B[3]), .B(B[2]), .ZN(n31) );
  XNOR2_X1 U32 ( .A(n54), .B(n64), .ZN(n52) );
  XOR2_X1 U33 ( .A(A[25]), .B(A[24]), .Z(n64) );
  XNOR2_X1 U48 ( .A(n52), .B(n65), .ZN(n50) );
  XNOR2_X1 U56 ( .A(n55), .B(n56), .ZN(n65) );
  XNOR2_X1 U57 ( .A(n66), .B(n34), .ZN(n1) );
  XNOR2_X1 U58 ( .A(n50), .B(n49), .ZN(n66) );
  XNOR2_X1 U59 ( .A(A[0]), .B(A[1]), .ZN(n54) );
endmodule


module NORGate_NX1_N32 ( A, B, Y );
  input [31:0] A;
  input [31:0] B;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21;

  OR3_X1 U1 ( .A1(n3), .A2(n1), .A3(n2), .ZN(n21) );
  NOR2_X1 U2 ( .A1(n4), .A2(n21), .ZN(Y) );
  NAND4_X1 U3 ( .A1(n5), .A2(n6), .A3(n7), .A4(n8), .ZN(n4) );
  NOR4_X1 U4 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n6) );
  NOR4_X1 U5 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n7) );
  NOR4_X1 U6 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n8) );
  NOR4_X1 U7 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n11) );
  NAND4_X1 U8 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .ZN(n3) );
  NOR4_X1 U9 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n12) );
  NOR4_X1 U10 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n9) );
  NOR4_X1 U11 ( .A1(A[30]), .A2(A[2]), .A3(A[29]), .A4(A[28]), .ZN(n10) );
  NAND4_X1 U12 ( .A1(n17), .A2(n18), .A3(n19), .A4(n20), .ZN(n1) );
  NAND4_X1 U13 ( .A1(n13), .A2(n14), .A3(n15), .A4(n16), .ZN(n2) );
  NOR4_X1 U14 ( .A1(B[12]), .A2(B[11]), .A3(B[10]), .A4(B[0]), .ZN(n13) );
  NOR4_X1 U15 ( .A1(B[16]), .A2(B[15]), .A3(B[14]), .A4(B[13]), .ZN(n14) );
  NOR4_X1 U16 ( .A1(B[1]), .A2(B[19]), .A3(B[18]), .A4(B[17]), .ZN(n15) );
  NOR4_X1 U17 ( .A1(B[23]), .A2(B[22]), .A3(B[21]), .A4(B[20]), .ZN(n16) );
  NOR4_X1 U18 ( .A1(B[9]), .A2(B[8]), .A3(B[7]), .A4(B[6]), .ZN(n20) );
  NOR4_X1 U19 ( .A1(B[5]), .A2(B[4]), .A3(B[3]), .A4(B[31]), .ZN(n19) );
  NOR4_X1 U20 ( .A1(B[30]), .A2(B[2]), .A3(B[29]), .A4(B[28]), .ZN(n18) );
  NOR4_X1 U21 ( .A1(B[27]), .A2(B[26]), .A3(B[25]), .A4(B[24]), .ZN(n17) );
  NOR4_X1 U22 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n5) );
endmodule


module Comparator_NBIT_DATA32 ( CMP_OpA, CMP_OpB, CMP_sgn_usgn, CMP_A_gt_B, 
        CMP_A_ge_B, CMP_A_lt_B, CMP_A_le_B, CMP_A_eq_B );
  input [31:0] CMP_OpA;
  input [31:0] CMP_OpB;
  input CMP_sgn_usgn;
  output CMP_A_gt_B, CMP_A_ge_B, CMP_A_lt_B, CMP_A_le_B, CMP_A_eq_B;
  wire   n325, s_en_mux, s_tmp_gt, s_tmp_lt, s_not_tmp_gt, s_not_tmp_lt, n44,
         n45, n46, n47, n48, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n81, n82, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n109, n110, n111, n112, n113, n114,
         n115, n116, n117, n118, n119, n120, n121, n122, n123, n124, n125,
         n126, n127, n128, n129, n130, n131, n132, n133, n134, n135, n136,
         n137, n138, n140, n141, n142, n143, n147, n148, n152, n153, n157,
         n158, n162, n163, n167, n168, n173, n174, n176, n178, n181, n182,
         n183, n184, n185, n139, n144, n145, n146, n149, n150, n151, n154,
         n155, n156, n159, n160, n161, n164, n165, n166, n169, n170, n171,
         n172, n175, n177, n179, n180, n186, n187, n188, n189, n190, n191,
         n192, n193, n194, n195, n196, n197, n198, n199, n200, n201, n202,
         n203, n204, n205, n206, n207, n208, n209, n210, n211, n212, n213,
         n214, n215, n216, n217, n218, n219, n220, n221, n222, n223, n224,
         n225, n226, n227, n228, n229, n230, n231, n232, n233, n234, n235,
         n236, n237, n238, n239, n240, n241, n242, n243, n244, n245, n246,
         n247, n248, n249, n250, n251, n252, n253, n254, n255, n256, n257,
         n258, n259, n260, n261, n262, n263, n264, n265, n266, n267, n268,
         n269, n270, n271, n272, n273, n274, n275, n276, n277, n278, n279,
         n280, n281, n282, n283, n284, n285, n286, n287, n288, n289, n290,
         n291, n292, n293, n294, n295, n296, n297, n298, n299, n300, n301,
         n302, n303, n304, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324;
  wire   [31:0] s_gt;
  wire   [31:0] s_lt;

  NAND3_X1 U185 ( .A1(n138), .A2(n213), .A3(CMP_OpB[0]), .ZN(n105) );
  XOR2_X1 U186 ( .A(CMP_OpB[1]), .B(CMP_OpA[1]), .Z(n140) );
  NAND3_X1 U203 ( .A1(n84), .A2(n168), .A3(n207), .ZN(n87) );
  NAND3_X1 U208 ( .A1(n74), .A2(n279), .A3(n204), .ZN(n176) );
  NAND3_X1 U209 ( .A1(n71), .A2(n178), .A3(n279), .ZN(n74) );
  NAND3_X1 U211 ( .A1(n68), .A2(n293), .A3(n205), .ZN(n181) );
  NAND3_X1 U212 ( .A1(n65), .A2(n183), .A3(n293), .ZN(n68) );
  ORGate_NX1_N32_2 OR_gt ( .A(s_gt), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .Y(s_tmp_gt) );
  ORGate_NX1_N32_1 OR_lt ( .A(s_lt), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .Y(s_tmp_lt) );
  Mux_1Bit_2X1_2 MUX_gt ( .port0(s_tmp_gt), .port1(s_not_tmp_gt), .sel(
        s_en_mux), .portY(n325) );
  Mux_1Bit_2X1_1 MUX_lt ( .port0(s_tmp_lt), .port1(s_not_tmp_lt), .sel(
        s_en_mux), .portY(CMP_A_lt_B) );
  NAND2_X1 U2 ( .A1(n75), .A2(n139), .ZN(n220) );
  AND2_X1 U3 ( .A1(n223), .A2(CMP_OpB[22]), .ZN(n139) );
  NAND2_X1 U4 ( .A1(n266), .A2(n287), .ZN(n144) );
  NAND2_X1 U5 ( .A1(n75), .A2(n145), .ZN(n78) );
  AND2_X1 U6 ( .A1(n223), .A2(CMP_OpB[22]), .ZN(n145) );
  NAND2_X1 U7 ( .A1(n149), .A2(n146), .ZN(n318) );
  INV_X32 U8 ( .A(n128), .ZN(n146) );
  AND3_X1 U9 ( .A1(n317), .A2(n207), .A3(n87), .ZN(n149) );
  AND2_X1 U10 ( .A1(n81), .A2(n288), .ZN(n150) );
  AND2_X1 U11 ( .A1(n81), .A2(n288), .ZN(n167) );
  NAND2_X1 U12 ( .A1(n141), .A2(CMP_OpA[2]), .ZN(n151) );
  AND2_X1 U13 ( .A1(n57), .A2(CMP_OpB[2]), .ZN(n154) );
  CLKBUF_X1 U14 ( .A(n57), .Z(n155) );
  AND2_X1 U15 ( .A1(CMP_OpB[1]), .A2(n140), .ZN(n156) );
  CLKBUF_X1 U16 ( .A(n238), .Z(n165) );
  CLKBUF_X1 U17 ( .A(n147), .Z(n297) );
  CLKBUF_X1 U18 ( .A(n228), .Z(n159) );
  CLKBUF_X1 U19 ( .A(n155), .Z(n160) );
  NAND3_X1 U20 ( .A1(n77), .A2(n173), .A3(n310), .ZN(n161) );
  AND2_X2 U21 ( .A1(n94), .A2(n196), .ZN(n157) );
  AND2_X2 U22 ( .A1(n100), .A2(n165), .ZN(n152) );
  NAND3_X1 U23 ( .A1(n65), .A2(n183), .A3(n293), .ZN(n164) );
  NAND2_X1 U24 ( .A1(n212), .A2(CMP_OpB[28]), .ZN(n166) );
  CLKBUF_X1 U25 ( .A(n132), .Z(n169) );
  NOR2_X1 U26 ( .A1(n302), .A2(n217), .ZN(n170) );
  NAND2_X1 U27 ( .A1(n184), .A2(CMP_OpA[29]), .ZN(n171) );
  XNOR2_X1 U28 ( .A(n172), .B(n175), .ZN(n48) );
  AND2_X1 U29 ( .A1(n147), .A2(CMP_OpA[7]), .ZN(n172) );
  AND2_X1 U30 ( .A1(n229), .A2(CMP_OpB[7]), .ZN(n175) );
  XNOR2_X1 U31 ( .A(n64), .B(n116), .ZN(n177) );
  XNOR2_X1 U32 ( .A(n263), .B(n231), .ZN(n179) );
  XNOR2_X1 U33 ( .A(n151), .B(n62), .ZN(n180) );
  AND2_X1 U34 ( .A1(n226), .A2(n289), .ZN(n244) );
  AND3_X1 U35 ( .A1(n99), .A2(n290), .A3(n315), .ZN(n238) );
  AND2_X1 U36 ( .A1(n290), .A2(n158), .ZN(n186) );
  AND2_X1 U37 ( .A1(n262), .A2(CMP_OpB[4]), .ZN(n187) );
  AND2_X1 U38 ( .A1(n244), .A2(n163), .ZN(n188) );
  CLKBUF_X1 U39 ( .A(n144), .Z(n189) );
  NAND2_X1 U40 ( .A1(n190), .A2(CMP_OpA[20]), .ZN(n309) );
  AND3_X1 U41 ( .A1(n161), .A2(n310), .A3(n228), .ZN(n190) );
  AND2_X1 U42 ( .A1(n75), .A2(n223), .ZN(n191) );
  AND2_X1 U43 ( .A1(n297), .A2(n148), .ZN(n192) );
  NAND2_X1 U44 ( .A1(n193), .A2(CMP_OpA[14]), .ZN(n319) );
  AND3_X1 U45 ( .A1(n93), .A2(n316), .A3(n244), .ZN(n193) );
  CLKBUF_X1 U46 ( .A(n111), .Z(n201) );
  NAND2_X1 U47 ( .A1(n229), .A2(CMP_OpB[7]), .ZN(n194) );
  BUF_X1 U48 ( .A(n237), .Z(n262) );
  AND3_X1 U49 ( .A1(n51), .A2(n297), .A3(n282), .ZN(n237) );
  AND3_X1 U50 ( .A1(n87), .A2(n317), .A3(n207), .ZN(n195) );
  CLKBUF_X1 U51 ( .A(n55), .Z(n224) );
  AND3_X1 U52 ( .A1(n93), .A2(n316), .A3(n244), .ZN(n196) );
  CLKBUF_X1 U53 ( .A(n319), .Z(n197) );
  AND2_X1 U54 ( .A1(CMP_OpA[1]), .A2(n140), .ZN(n198) );
  NAND3_X1 U55 ( .A1(n138), .A2(n213), .A3(CMP_OpB[0]), .ZN(n199) );
  NAND2_X1 U56 ( .A1(n147), .A2(CMP_OpA[7]), .ZN(n200) );
  CLKBUF_X1 U57 ( .A(n164), .Z(n202) );
  CLKBUF_X1 U58 ( .A(n74), .Z(n203) );
  XNOR2_X1 U59 ( .A(n72), .B(n120), .ZN(n204) );
  XNOR2_X1 U60 ( .A(n166), .B(n117), .ZN(n205) );
  CLKBUF_X1 U61 ( .A(n307), .Z(n206) );
  CLKBUF_X1 U62 ( .A(n150), .Z(n207) );
  CLKBUF_X1 U63 ( .A(n166), .Z(n208) );
  AND2_X1 U64 ( .A1(n262), .A2(CMP_OpA[4]), .ZN(n209) );
  CLKBUF_X1 U65 ( .A(n47), .Z(n210) );
  CLKBUF_X1 U66 ( .A(n323), .Z(n211) );
  AND2_X1 U67 ( .A1(n177), .A2(n243), .ZN(n212) );
  AND2_X1 U68 ( .A1(n61), .A2(n296), .ZN(n213) );
  NAND2_X1 U69 ( .A1(n214), .A2(CMP_OpA[11]), .ZN(n323) );
  AND3_X1 U70 ( .A1(n99), .A2(n290), .A3(n315), .ZN(n214) );
  XNOR2_X1 U71 ( .A(n250), .B(n222), .ZN(n215) );
  XNOR2_X1 U72 ( .A(n267), .B(n256), .ZN(n216) );
  XNOR2_X1 U73 ( .A(CMP_OpA[30]), .B(n60), .ZN(n217) );
  NAND2_X1 U74 ( .A1(n218), .A2(CMP_OpA[8]), .ZN(n324) );
  AND3_X1 U75 ( .A1(n45), .A2(n299), .A3(n307), .ZN(n218) );
  CLKBUF_X1 U76 ( .A(n157), .Z(n290) );
  AND2_X1 U77 ( .A1(n180), .A2(n296), .ZN(n303) );
  NAND3_X1 U78 ( .A1(n77), .A2(n173), .A3(n310), .ZN(n219) );
  CLKBUF_X1 U79 ( .A(n87), .Z(n221) );
  CLKBUF_X1 U80 ( .A(n103), .Z(n222) );
  CLKBUF_X1 U81 ( .A(n174), .Z(n223) );
  NAND2_X1 U82 ( .A1(CMP_OpB[23]), .A2(n174), .ZN(n225) );
  XNOR2_X1 U83 ( .A(n89), .B(n318), .ZN(n226) );
  CLKBUF_X1 U84 ( .A(n48), .Z(n227) );
  XNOR2_X1 U85 ( .A(n220), .B(n144), .ZN(n228) );
  AND2_X1 U86 ( .A1(n46), .A2(n252), .ZN(n229) );
  BUF_X1 U87 ( .A(n195), .Z(n289) );
  NAND2_X1 U88 ( .A1(n180), .A2(n230), .ZN(n138) );
  AND2_X1 U89 ( .A1(n296), .A2(n140), .ZN(n230) );
  NAND2_X1 U90 ( .A1(n237), .A2(CMP_OpA[5]), .ZN(n231) );
  CLKBUF_X1 U91 ( .A(n200), .Z(n232) );
  AND2_X1 U92 ( .A1(n303), .A2(n140), .ZN(n233) );
  CLKBUF_X1 U93 ( .A(n64), .Z(n234) );
  NAND2_X1 U94 ( .A1(n289), .A2(CMP_OpB[17]), .ZN(n235) );
  CLKBUF_X1 U95 ( .A(CMP_OpA[31]), .Z(n236) );
  AND2_X1 U96 ( .A1(n46), .A2(n252), .ZN(n147) );
  AND3_X1 U97 ( .A1(n45), .A2(n299), .A3(n307), .ZN(n239) );
  NAND2_X1 U98 ( .A1(n240), .A2(CMP_OpA[5]), .ZN(n320) );
  AND3_X1 U99 ( .A1(n51), .A2(n297), .A3(n282), .ZN(n240) );
  CLKBUF_X1 U100 ( .A(n120), .Z(n241) );
  CLKBUF_X1 U101 ( .A(n317), .Z(n242) );
  NOR2_X1 U102 ( .A1(n114), .A2(n58), .ZN(n243) );
  CLKBUF_X1 U103 ( .A(n117), .Z(n245) );
  CLKBUF_X1 U104 ( .A(n161), .Z(n246) );
  AND2_X1 U105 ( .A1(n88), .A2(n289), .ZN(n162) );
  AND3_X1 U106 ( .A1(n219), .A2(n310), .A3(n228), .ZN(n247) );
  CLKBUF_X1 U107 ( .A(n324), .Z(n248) );
  NAND2_X1 U108 ( .A1(n296), .A2(CMP_OpB[2]), .ZN(n249) );
  CLKBUF_X1 U109 ( .A(n135), .Z(n250) );
  CLKBUF_X1 U110 ( .A(n82), .Z(n251) );
  CLKBUF_X1 U111 ( .A(n239), .Z(n252) );
  NAND2_X1 U112 ( .A1(n227), .A2(n192), .ZN(n253) );
  CLKBUF_X1 U113 ( .A(n99), .Z(n254) );
  CLKBUF_X1 U114 ( .A(n249), .Z(n255) );
  XNOR2_X1 U115 ( .A(n91), .B(n256), .ZN(n316) );
  NAND2_X1 U116 ( .A1(CMP_OpA[16]), .A2(n244), .ZN(n256) );
  CLKBUF_X1 U117 ( .A(n126), .Z(n257) );
  CLKBUF_X1 U118 ( .A(n93), .Z(n258) );
  NAND2_X1 U119 ( .A1(n165), .A2(CMP_OpB[11]), .ZN(n259) );
  AND3_X1 U120 ( .A1(n164), .A2(n293), .A3(n205), .ZN(n260) );
  CLKBUF_X1 U121 ( .A(n171), .Z(n261) );
  NAND2_X1 U122 ( .A1(n52), .A2(n209), .ZN(n111) );
  NAND2_X1 U123 ( .A1(n237), .A2(CMP_OpB[5]), .ZN(n263) );
  CLKBUF_X1 U124 ( .A(n97), .Z(n264) );
  NOR2_X1 U125 ( .A1(n199), .A2(n137), .ZN(n265) );
  NAND2_X1 U126 ( .A1(n52), .A2(n187), .ZN(n55) );
  XNOR2_X1 U127 ( .A(n322), .B(n225), .ZN(n266) );
  OR2_X2 U128 ( .A1(n304), .A2(n181), .ZN(n70) );
  CLKBUF_X1 U129 ( .A(n91), .Z(n267) );
  NAND2_X1 U130 ( .A1(CMP_OpB[8]), .A2(n252), .ZN(n268) );
  NAND2_X1 U131 ( .A1(CMP_OpA[2]), .A2(n296), .ZN(n269) );
  CLKBUF_X1 U132 ( .A(n114), .Z(n270) );
  XNOR2_X1 U133 ( .A(n224), .B(n201), .ZN(n271) );
  CLKBUF_X1 U134 ( .A(n95), .Z(n272) );
  XNOR2_X1 U135 ( .A(n263), .B(n231), .ZN(n273) );
  XNOR2_X1 U136 ( .A(n70), .B(n280), .ZN(n274) );
  XNOR2_X1 U137 ( .A(n211), .B(n259), .ZN(n275) );
  XNOR2_X1 U138 ( .A(n269), .B(n249), .ZN(n276) );
  CLKBUF_X1 U139 ( .A(n226), .Z(n277) );
  XNOR2_X1 U140 ( .A(n320), .B(n53), .ZN(n52) );
  CLKBUF_X1 U141 ( .A(n177), .Z(n278) );
  AND2_X1 U142 ( .A1(n283), .A2(n260), .ZN(n279) );
  INV_X1 U143 ( .A(CMP_OpA[3]), .ZN(n112) );
  INV_X1 U144 ( .A(CMP_OpA[26]), .ZN(n119) );
  AND2_X1 U145 ( .A1(n303), .A2(n198), .ZN(s_gt[1]) );
  INV_X1 U146 ( .A(CMP_OpA[6]), .ZN(n109) );
  INV_X1 U147 ( .A(CMP_OpA[21]), .ZN(n124) );
  INV_X1 U148 ( .A(CMP_OpA[18]), .ZN(n127) );
  INV_X1 U149 ( .A(CMP_OpA[15]), .ZN(n130) );
  INV_X1 U150 ( .A(CMP_OpA[12]), .ZN(n133) );
  INV_X1 U151 ( .A(CMP_OpA[17]), .ZN(n128) );
  INV_X1 U152 ( .A(CMP_OpA[11]), .ZN(n134) );
  INV_X1 U153 ( .A(CMP_OpA[23]), .ZN(n122) );
  INV_X1 U154 ( .A(CMP_OpA[20]), .ZN(n125) );
  INV_X1 U155 ( .A(CMP_OpA[14]), .ZN(n131) );
  INV_X1 U156 ( .A(CMP_OpA[24]), .ZN(n121) );
  INV_X1 U157 ( .A(CMP_OpA[5]), .ZN(n110) );
  INV_X1 U158 ( .A(CMP_OpA[8]), .ZN(n107) );
  INV_X1 U159 ( .A(CMP_OpA[0]), .ZN(n137) );
  INV_X1 U160 ( .A(CMP_OpA[27]), .ZN(n118) );
  INV_X1 U161 ( .A(CMP_OpA[9]), .ZN(n106) );
  XNOR2_X1 U162 ( .A(n70), .B(n280), .ZN(n69) );
  OR2_X1 U163 ( .A1(n181), .A2(n119), .ZN(n280) );
  XNOR2_X1 U164 ( .A(n89), .B(n318), .ZN(n88) );
  XNOR2_X1 U165 ( .A(n73), .B(CMP_OpA[24]), .ZN(n178) );
  XNOR2_X1 U166 ( .A(n79), .B(CMP_OpA[21]), .ZN(n173) );
  XNOR2_X1 U167 ( .A(n86), .B(CMP_OpA[18]), .ZN(n168) );
  XNOR2_X1 U168 ( .A(n67), .B(CMP_OpA[27]), .ZN(n183) );
  XNOR2_X1 U169 ( .A(n56), .B(CMP_OpA[3]), .ZN(n143) );
  AND2_X1 U170 ( .A1(n299), .A2(n153), .ZN(n281) );
  INV_X1 U171 ( .A(CMP_OpB[31]), .ZN(n321) );
  INV_X1 U172 ( .A(CMP_OpB[26]), .ZN(n304) );
  AND2_X1 U173 ( .A1(n303), .A2(n156), .ZN(s_lt[1]) );
  INV_X1 U174 ( .A(CMP_OpB[27]), .ZN(n67) );
  INV_X1 U175 ( .A(CMP_OpB[21]), .ZN(n79) );
  INV_X1 U176 ( .A(CMP_OpB[24]), .ZN(n73) );
  INV_X1 U177 ( .A(CMP_OpB[18]), .ZN(n86) );
  INV_X1 U178 ( .A(CMP_OpB[30]), .ZN(n60) );
  INV_X1 U179 ( .A(CMP_OpB[15]), .ZN(n92) );
  INV_X1 U180 ( .A(CMP_OpB[12]), .ZN(n98) );
  INV_X1 U181 ( .A(CMP_OpB[6]), .ZN(n50) );
  INV_X1 U182 ( .A(CMP_OpB[9]), .ZN(n44) );
  INV_X1 U183 ( .A(CMP_OpB[3]), .ZN(n56) );
  XNOR2_X1 U184 ( .A(n72), .B(n120), .ZN(n71) );
  XNOR2_X1 U187 ( .A(n200), .B(n194), .ZN(n282) );
  CLKBUF_X1 U188 ( .A(n274), .Z(n283) );
  AND2_X1 U189 ( .A1(CMP_OpB[25]), .A2(n260), .ZN(n284) );
  AND2_X1 U190 ( .A1(CMP_OpA[25]), .A2(n260), .ZN(n285) );
  CLKBUF_X1 U191 ( .A(n220), .Z(n286) );
  AND2_X1 U192 ( .A1(CMP_OpA[22]), .A2(n223), .ZN(n287) );
  CLKBUF_X1 U193 ( .A(n247), .Z(n288) );
  CLKBUF_X1 U194 ( .A(n191), .Z(n310) );
  XNOR2_X1 U195 ( .A(n272), .B(n197), .ZN(n291) );
  XNOR2_X1 U196 ( .A(n95), .B(n319), .ZN(n94) );
  CLKBUF_X1 U197 ( .A(n212), .Z(n293) );
  XNOR2_X1 U198 ( .A(n64), .B(n171), .ZN(n63) );
  CLKBUF_X1 U199 ( .A(n70), .Z(n292) );
  AND2_X1 U200 ( .A1(n63), .A2(n243), .ZN(n182) );
  CLKBUF_X1 U201 ( .A(n194), .Z(n294) );
  CLKBUF_X1 U202 ( .A(n72), .Z(n295) );
  AND2_X1 U204 ( .A1(n57), .A2(n142), .ZN(n296) );
  AND2_X1 U205 ( .A1(n57), .A2(n142), .ZN(n141) );
  CLKBUF_X1 U206 ( .A(n152), .Z(n299) );
  AND2_X1 U207 ( .A1(n143), .A2(n311), .ZN(n298) );
  INV_X1 U210 ( .A(n303), .ZN(n136) );
  CLKBUF_X1 U213 ( .A(n225), .Z(n300) );
  NAND2_X1 U214 ( .A1(n215), .A2(n281), .ZN(n301) );
  XNOR2_X1 U215 ( .A(CMP_OpA[31]), .B(n321), .ZN(n302) );
  NAND2_X1 U216 ( .A1(n274), .A2(n284), .ZN(n72) );
  NAND2_X1 U217 ( .A1(n69), .A2(n285), .ZN(n120) );
  NAND2_X1 U218 ( .A1(n141), .A2(CMP_OpA[2]), .ZN(n115) );
  NAND2_X1 U219 ( .A1(n154), .A2(n142), .ZN(n62) );
  XNOR2_X1 U220 ( .A(n115), .B(n62), .ZN(n61) );
  NAND2_X1 U221 ( .A1(CMP_A_lt_B), .A2(n185), .ZN(CMP_A_ge_B) );
  INV_X1 U222 ( .A(s_tmp_lt), .ZN(s_not_tmp_lt) );
  INV_X1 U223 ( .A(CMP_OpA[30]), .ZN(n113) );
  CLKBUF_X1 U224 ( .A(n325), .Z(CMP_A_gt_B) );
  NAND2_X1 U225 ( .A1(n48), .A2(n192), .ZN(n51) );
  NAND2_X1 U226 ( .A1(n102), .A2(n281), .ZN(n45) );
  CLKBUF_X1 U227 ( .A(n302), .Z(n306) );
  XNOR2_X1 U228 ( .A(n103), .B(n135), .ZN(n307) );
  XNOR2_X1 U229 ( .A(n50), .B(CMP_OpA[6]), .ZN(n148) );
  XNOR2_X1 U230 ( .A(n44), .B(CMP_OpA[9]), .ZN(n153) );
  INV_X1 U231 ( .A(s_tmp_gt), .ZN(s_not_tmp_gt) );
  NOR2_X1 U232 ( .A1(CMP_A_lt_B), .A2(CMP_A_gt_B), .ZN(CMP_A_eq_B) );
  INV_X1 U233 ( .A(n325), .ZN(n185) );
  INV_X1 U234 ( .A(n270), .ZN(n59) );
  OR2_X1 U235 ( .A1(n185), .A2(CMP_A_lt_B), .ZN(CMP_A_le_B) );
  XNOR2_X1 U236 ( .A(n135), .B(n103), .ZN(n102) );
  INV_X1 U237 ( .A(n176), .ZN(n174) );
  CLKBUF_X1 U238 ( .A(n81), .Z(n308) );
  XNOR2_X1 U239 ( .A(n82), .B(n309), .ZN(n81) );
  NAND2_X1 U240 ( .A1(n157), .A2(CMP_OpB[13]), .ZN(n97) );
  NAND2_X1 U241 ( .A1(n152), .A2(CMP_OpA[10]), .ZN(n135) );
  NAND2_X1 U242 ( .A1(n152), .A2(CMP_OpB[10]), .ZN(n103) );
  NOR2_X1 U243 ( .A1(n44), .A2(n301), .ZN(s_lt[9]) );
  NOR2_X1 U244 ( .A1(n206), .A2(n222), .ZN(s_lt[10]) );
  NOR2_X1 U245 ( .A1(n50), .A2(n253), .ZN(s_lt[6]) );
  NOR2_X1 U246 ( .A1(n106), .A2(n301), .ZN(s_gt[9]) );
  NOR2_X1 U247 ( .A1(n109), .A2(n253), .ZN(s_gt[6]) );
  AND2_X1 U248 ( .A1(n273), .A2(n262), .ZN(n311) );
  AND2_X1 U249 ( .A1(n54), .A2(n311), .ZN(n142) );
  NAND2_X1 U250 ( .A1(n96), .A2(n186), .ZN(n99) );
  NAND2_X1 U251 ( .A1(n90), .A2(n188), .ZN(n93) );
  NOR2_X1 U252 ( .A1(n114), .A2(n58), .ZN(n312) );
  XNOR2_X1 U253 ( .A(n268), .B(n248), .ZN(n313) );
  CLKBUF_X1 U254 ( .A(n266), .Z(n314) );
  XNOR2_X1 U255 ( .A(n97), .B(n132), .ZN(n315) );
  BUF_X1 U256 ( .A(n84), .Z(n317) );
  XNOR2_X1 U257 ( .A(n98), .B(CMP_OpA[12]), .ZN(n158) );
  XNOR2_X1 U258 ( .A(n92), .B(CMP_OpA[15]), .ZN(n163) );
  XNOR2_X1 U259 ( .A(n66), .B(n117), .ZN(n65) );
  NOR2_X1 U260 ( .A1(n307), .A2(n250), .ZN(s_gt[10]) );
  XNOR2_X1 U261 ( .A(CMP_OpA[31]), .B(n321), .ZN(n58) );
  XNOR2_X1 U262 ( .A(n76), .B(n322), .ZN(n75) );
  OR2_X1 U263 ( .A1(n176), .A2(n122), .ZN(n322) );
  XNOR2_X1 U264 ( .A(n323), .B(n101), .ZN(n100) );
  XNOR2_X1 U265 ( .A(n47), .B(n324), .ZN(n46) );
  NOR2_X1 U266 ( .A1(n179), .A2(n263), .ZN(s_lt[5]) );
  NOR2_X1 U267 ( .A1(n283), .A2(n292), .ZN(s_lt[26]) );
  NOR2_X1 U268 ( .A1(n73), .A2(n203), .ZN(s_lt[24]) );
  NOR2_X1 U269 ( .A1(n56), .A2(n160), .ZN(s_lt[3]) );
  NOR2_X1 U270 ( .A1(n282), .A2(n294), .ZN(s_lt[7]) );
  NOR2_X1 U271 ( .A1(n179), .A2(n110), .ZN(s_gt[5]) );
  NOR2_X1 U272 ( .A1(n119), .A2(n283), .ZN(s_gt[26]) );
  NOR2_X1 U273 ( .A1(n121), .A2(n203), .ZN(s_gt[24]) );
  NOR2_X1 U274 ( .A1(n112), .A2(n155), .ZN(s_gt[3]) );
  NOR2_X1 U275 ( .A1(n282), .A2(n232), .ZN(s_gt[7]) );
  NAND2_X1 U276 ( .A1(n157), .A2(CMP_OpA[13]), .ZN(n132) );
  NAND2_X1 U277 ( .A1(n162), .A2(CMP_OpB[16]), .ZN(n91) );
  NAND2_X1 U278 ( .A1(n212), .A2(CMP_OpB[28]), .ZN(n66) );
  XNOR2_X1 U279 ( .A(n91), .B(n129), .ZN(n90) );
  NAND2_X1 U280 ( .A1(n162), .A2(CMP_OpA[16]), .ZN(n129) );
  XNOR2_X1 U281 ( .A(n123), .B(n78), .ZN(n77) );
  NAND2_X1 U282 ( .A1(n266), .A2(n287), .ZN(n123) );
  NAND2_X1 U283 ( .A1(n182), .A2(CMP_OpA[28]), .ZN(n117) );
  XNOR2_X1 U284 ( .A(n85), .B(n126), .ZN(n84) );
  NAND2_X1 U285 ( .A1(CMP_OpB[19]), .A2(n150), .ZN(n85) );
  XNOR2_X1 U286 ( .A(CMP_OpA[30]), .B(n60), .ZN(n114) );
  NAND2_X1 U287 ( .A1(n238), .A2(CMP_OpB[11]), .ZN(n101) );
  AND2_X1 U288 ( .A1(CMP_sgn_usgn), .A2(n306), .ZN(s_en_mux) );
  NOR3_X1 U289 ( .A1(n306), .A2(n59), .A3(n60), .ZN(s_lt[30]) );
  NOR2_X1 U290 ( .A1(n98), .A2(n254), .ZN(s_lt[12]) );
  NOR2_X1 U291 ( .A1(n314), .A2(n300), .ZN(s_lt[23]) );
  NOR2_X1 U292 ( .A1(n92), .A2(n258), .ZN(s_lt[15]) );
  NOR2_X1 U293 ( .A1(n133), .A2(n254), .ZN(s_gt[12]) );
  NOR2_X1 U294 ( .A1(n314), .A2(n122), .ZN(s_gt[23]) );
  NOR3_X1 U295 ( .A1(n306), .A2(n59), .A3(n113), .ZN(s_gt[30]) );
  NOR2_X1 U296 ( .A1(n79), .A2(n246), .ZN(s_lt[21]) );
  AND2_X1 U297 ( .A1(n306), .A2(CMP_OpB[31]), .ZN(s_lt[31]) );
  NOR2_X1 U298 ( .A1(n130), .A2(n258), .ZN(s_gt[15]) );
  NOR2_X1 U299 ( .A1(n271), .A2(n201), .ZN(s_gt[4]) );
  NOR2_X1 U300 ( .A1(n124), .A2(n246), .ZN(s_gt[21]) );
  NAND2_X1 U301 ( .A1(n54), .A2(n298), .ZN(n57) );
  NOR2_X1 U302 ( .A1(n302), .A2(n217), .ZN(n184) );
  NOR2_X1 U303 ( .A1(n67), .A2(n202), .ZN(s_lt[27]) );
  NOR2_X1 U304 ( .A1(n204), .A2(n295), .ZN(s_lt[25]) );
  NOR2_X1 U305 ( .A1(n118), .A2(n202), .ZN(s_gt[27]) );
  NOR2_X1 U306 ( .A1(n242), .A2(n85), .ZN(s_lt[19]) );
  NOR2_X1 U307 ( .A1(n86), .A2(n221), .ZN(s_lt[18]) );
  NOR2_X1 U308 ( .A1(n277), .A2(n235), .ZN(s_lt[17]) );
  NOR2_X1 U309 ( .A1(n308), .A2(n251), .ZN(s_lt[20]) );
  NOR2_X1 U310 ( .A1(n242), .A2(n257), .ZN(s_gt[19]) );
  NOR2_X1 U311 ( .A1(n204), .A2(n241), .ZN(s_gt[25]) );
  NOR2_X1 U312 ( .A1(n127), .A2(n221), .ZN(s_gt[18]) );
  NOR2_X1 U313 ( .A1(n308), .A2(n125), .ZN(s_gt[20]) );
  NOR2_X1 U314 ( .A1(n277), .A2(n128), .ZN(s_gt[17]) );
  NOR2_X1 U315 ( .A1(n105), .A2(n137), .ZN(n104) );
  NAND2_X1 U316 ( .A1(n312), .A2(CMP_OpB[29]), .ZN(n64) );
  NAND2_X1 U317 ( .A1(n170), .A2(CMP_OpA[29]), .ZN(n116) );
  XNOR2_X1 U318 ( .A(n132), .B(n97), .ZN(n96) );
  NAND2_X1 U319 ( .A1(n167), .A2(CMP_OpA[19]), .ZN(n126) );
  NAND2_X1 U320 ( .A1(n239), .A2(CMP_OpB[8]), .ZN(n47) );
  NAND2_X1 U321 ( .A1(n196), .A2(CMP_OpB[14]), .ZN(n95) );
  NAND2_X1 U322 ( .A1(n195), .A2(CMP_OpB[17]), .ZN(n89) );
  NAND2_X1 U323 ( .A1(n247), .A2(CMP_OpB[20]), .ZN(n82) );
  NAND2_X1 U324 ( .A1(n174), .A2(CMP_OpB[23]), .ZN(n76) );
  NAND2_X1 U325 ( .A1(n240), .A2(CMP_OpB[5]), .ZN(n53) );
  NOR2_X1 U326 ( .A1(n216), .A2(n267), .ZN(s_lt[16]) );
  NOR2_X1 U327 ( .A1(n276), .A2(n255), .ZN(s_lt[2]) );
  NOR2_X1 U328 ( .A1(n271), .A2(n224), .ZN(s_lt[4]) );
  NOR2_X1 U329 ( .A1(n313), .A2(n210), .ZN(s_lt[8]) );
  NOR2_X1 U330 ( .A1(n278), .A2(n234), .ZN(s_lt[29]) );
  NOR2_X1 U331 ( .A1(n275), .A2(n259), .ZN(s_lt[11]) );
  NOR2_X1 U332 ( .A1(n205), .A2(n208), .ZN(s_lt[28]) );
  NOR2_X1 U333 ( .A1(n159), .A2(n286), .ZN(s_lt[22]) );
  NOR2_X1 U334 ( .A1(n265), .A2(n199), .ZN(s_lt[0]) );
  NOR2_X1 U335 ( .A1(n291), .A2(n272), .ZN(s_lt[14]) );
  NOR2_X1 U336 ( .A1(n264), .A2(n315), .ZN(s_lt[13]) );
  NOR2_X1 U337 ( .A1(n216), .A2(n129), .ZN(s_gt[16]) );
  NOR2_X1 U338 ( .A1(n276), .A2(n269), .ZN(s_gt[2]) );
  NOR2_X1 U339 ( .A1(n313), .A2(n107), .ZN(s_gt[8]) );
  NOR2_X1 U340 ( .A1(n278), .A2(n261), .ZN(s_gt[29]) );
  NOR2_X1 U341 ( .A1(n275), .A2(n134), .ZN(s_gt[11]) );
  NOR2_X1 U342 ( .A1(n205), .A2(n245), .ZN(s_gt[28]) );
  NOR2_X1 U343 ( .A1(n159), .A2(n189), .ZN(s_gt[22]) );
  NOR4_X1 U344 ( .A1(n104), .A2(n233), .A3(n136), .A4(n137), .ZN(s_gt[0]) );
  NOR2_X1 U345 ( .A1(n291), .A2(n131), .ZN(s_gt[14]) );
  NOR2_X1 U346 ( .A1(n315), .A2(n169), .ZN(s_gt[13]) );
  AND2_X1 U347 ( .A1(n306), .A2(n236), .ZN(s_gt[31]) );
  XNOR2_X1 U348 ( .A(n55), .B(n111), .ZN(n54) );
endmodule


module CarrySelect_N32_K4 ( A, B, Cin, S );
  input [31:0] A;
  input [31:0] B;
  input [7:0] Cin;
  output [31:0] S;


  CarrySelectBlock_N4_0 CSB_i_0 ( .A(A[3:0]), .B(B[3:0]), .Cin(Cin[0]), .S(
        S[3:0]) );
  CarrySelectBlock_N4_7 CSB_i_4 ( .A(A[7:4]), .B(B[7:4]), .Cin(Cin[1]), .S(
        S[7:4]) );
  CarrySelectBlock_N4_6 CSB_i_8 ( .A(A[11:8]), .B(B[11:8]), .Cin(Cin[2]), .S(
        S[11:8]) );
  CarrySelectBlock_N4_5 CSB_i_12 ( .A(A[15:12]), .B(B[15:12]), .Cin(Cin[3]), 
        .S(S[15:12]) );
  CarrySelectBlock_N4_4 CSB_i_16 ( .A(A[19:16]), .B(B[19:16]), .Cin(Cin[4]), 
        .S(S[19:16]) );
  CarrySelectBlock_N4_3 CSB_i_20 ( .A(A[23:20]), .B(B[23:20]), .Cin(Cin[5]), 
        .S(S[23:20]) );
  CarrySelectBlock_N4_2 CSB_i_24 ( .A(A[27:24]), .B(B[27:24]), .Cin(Cin[6]), 
        .S(S[27:24]) );
  CarrySelectBlock_N4_1 CSB_i_28 ( .A(A[31:28]), .B(B[31:28]), .Cin(Cin[7]), 
        .S(S[31:28]) );
endmodule


module CarryGenerator_N32_K8 ( A, B, c_in, CarryVector );
  input [31:0] A;
  input [31:0] B;
  output [7:0] CarryVector;
  input c_in;
  wire   \P_mat[1][32] , \P_mat[1][31] , \P_mat[1][30] , \P_mat[1][29] ,
         \P_mat[1][28] , \P_mat[1][27] , \P_mat[1][26] , \P_mat[1][25] ,
         \P_mat[1][24] , \P_mat[1][23] , \P_mat[1][22] , \P_mat[1][21] ,
         \P_mat[1][20] , \P_mat[1][19] , \P_mat[1][18] , \P_mat[1][17] ,
         \P_mat[1][16] , \P_mat[1][15] , \P_mat[1][14] , \P_mat[1][13] ,
         \P_mat[1][12] , \P_mat[1][11] , \P_mat[1][10] , \P_mat[1][9] ,
         \P_mat[1][8] , \P_mat[1][7] , \P_mat[1][6] , \P_mat[1][5] ,
         \P_mat[1][4] , \P_mat[1][3] , \P_mat[1][2] , \P_mat[2][32] ,
         \P_mat[2][30] , \P_mat[2][28] , \P_mat[2][26] , \P_mat[2][24] ,
         \P_mat[2][22] , \P_mat[2][20] , \P_mat[2][18] , \P_mat[2][16] ,
         \P_mat[2][14] , \P_mat[2][12] , \P_mat[2][10] , \P_mat[2][8] ,
         \P_mat[2][6] , \P_mat[2][4] , \P_mat[3][32] , \P_mat[3][28] ,
         \P_mat[3][24] , \P_mat[3][20] , \P_mat[3][16] , \P_mat[3][12] ,
         \P_mat[3][8] , \P_mat[4][32] , \P_mat[4][24] , \P_mat[4][16] ,
         \P_mat[5][32] , \P_mat[5][28] , \G_mat[1][32] , \G_mat[1][31] ,
         \G_mat[1][30] , \G_mat[1][29] , \G_mat[1][28] , \G_mat[1][27] ,
         \G_mat[1][26] , \G_mat[1][25] , \G_mat[1][24] , \G_mat[1][23] ,
         \G_mat[1][22] , \G_mat[1][21] , \G_mat[1][20] , \G_mat[1][19] ,
         \G_mat[1][18] , \G_mat[1][17] , \G_mat[1][16] , \G_mat[1][15] ,
         \G_mat[1][14] , \G_mat[1][13] , \G_mat[1][12] , \G_mat[1][11] ,
         \G_mat[1][10] , \G_mat[1][9] , \G_mat[1][8] , \G_mat[1][7] ,
         \G_mat[1][6] , \G_mat[1][5] , \G_mat[1][4] , \G_mat[1][3] ,
         \G_mat[1][2] , \G_mat[1][1] , \G_mat[2][32] , \G_mat[2][30] ,
         \G_mat[2][28] , \G_mat[2][26] , \G_mat[2][24] , \G_mat[2][22] ,
         \G_mat[2][20] , \G_mat[2][18] , \G_mat[2][16] , \G_mat[2][14] ,
         \G_mat[2][12] , \G_mat[2][10] , \G_mat[2][8] , \G_mat[2][6] ,
         \G_mat[2][4] , \G_mat[2][2] , \G_mat[3][32] , \G_mat[3][28] ,
         \G_mat[3][24] , \G_mat[3][20] , \G_mat[3][16] , \G_mat[3][12] ,
         \G_mat[3][8] , \G_mat[4][32] , \G_mat[4][24] , \G_mat[4][16] ,
         \G_mat[5][32] , \G_mat[5][28] ;
  wire   SYNOPSYS_UNCONNECTED__0;

  PG_network_N32_1 PG_net ( .A(A), .B(B), .c_in(c_in), .G({\G_mat[1][32] , 
        \G_mat[1][31] , \G_mat[1][30] , \G_mat[1][29] , \G_mat[1][28] , 
        \G_mat[1][27] , \G_mat[1][26] , \G_mat[1][25] , \G_mat[1][24] , 
        \G_mat[1][23] , \G_mat[1][22] , \G_mat[1][21] , \G_mat[1][20] , 
        \G_mat[1][19] , \G_mat[1][18] , \G_mat[1][17] , \G_mat[1][16] , 
        \G_mat[1][15] , \G_mat[1][14] , \G_mat[1][13] , \G_mat[1][12] , 
        \G_mat[1][11] , \G_mat[1][10] , \G_mat[1][9] , \G_mat[1][8] , 
        \G_mat[1][7] , \G_mat[1][6] , \G_mat[1][5] , \G_mat[1][4] , 
        \G_mat[1][3] , \G_mat[1][2] , \G_mat[1][1] }), .P({\P_mat[1][32] , 
        \P_mat[1][31] , \P_mat[1][30] , \P_mat[1][29] , \P_mat[1][28] , 
        \P_mat[1][27] , \P_mat[1][26] , \P_mat[1][25] , \P_mat[1][24] , 
        \P_mat[1][23] , \P_mat[1][22] , \P_mat[1][21] , \P_mat[1][20] , 
        \P_mat[1][19] , \P_mat[1][18] , \P_mat[1][17] , \P_mat[1][16] , 
        \P_mat[1][15] , \P_mat[1][14] , \P_mat[1][13] , \P_mat[1][12] , 
        \P_mat[1][11] , \P_mat[1][10] , \P_mat[1][9] , \P_mat[1][8] , 
        \P_mat[1][7] , \P_mat[1][6] , \P_mat[1][5] , \P_mat[1][4] , 
        \P_mat[1][3] , \P_mat[1][2] , SYNOPSYS_UNCONNECTED__0}) );
  GeneralGenerate_10 PM0_1_1 ( .G_ik(\G_mat[1][2] ), .P_ik(\P_mat[1][2] ), 
        .G_km1_j(\G_mat[1][1] ), .G_ij(\G_mat[2][2] ) );
  GeneralPropagate_0 PM2_1_2 ( .G_ik(\G_mat[1][4] ), .P_ik(\P_mat[1][4] ), 
        .G_km1_j(\G_mat[1][3] ), .P_km1_j(\P_mat[1][3] ), .G_ij(\G_mat[2][4] ), 
        .P_ij(\P_mat[2][4] ) );
  GeneralPropagate_26 PM2_1_3 ( .G_ik(\G_mat[1][6] ), .P_ik(\P_mat[1][6] ), 
        .G_km1_j(\G_mat[1][5] ), .P_km1_j(\P_mat[1][5] ), .G_ij(\G_mat[2][6] ), 
        .P_ij(\P_mat[2][6] ) );
  GeneralPropagate_25 PM2_1_4 ( .G_ik(\G_mat[1][8] ), .P_ik(\P_mat[1][8] ), 
        .G_km1_j(\G_mat[1][7] ), .P_km1_j(\P_mat[1][7] ), .G_ij(\G_mat[2][8] ), 
        .P_ij(\P_mat[2][8] ) );
  GeneralPropagate_24 PM2_1_5 ( .G_ik(\G_mat[1][10] ), .P_ik(\P_mat[1][10] ), 
        .G_km1_j(\G_mat[1][9] ), .P_km1_j(\P_mat[1][9] ), .G_ij(\G_mat[2][10] ), .P_ij(\P_mat[2][10] ) );
  GeneralPropagate_23 PM2_1_6 ( .G_ik(\G_mat[1][12] ), .P_ik(\P_mat[1][12] ), 
        .G_km1_j(\G_mat[1][11] ), .P_km1_j(\P_mat[1][11] ), .G_ij(
        \G_mat[2][12] ), .P_ij(\P_mat[2][12] ) );
  GeneralPropagate_22 PM2_1_7 ( .G_ik(\G_mat[1][14] ), .P_ik(\P_mat[1][14] ), 
        .G_km1_j(\G_mat[1][13] ), .P_km1_j(\P_mat[1][13] ), .G_ij(
        \G_mat[2][14] ), .P_ij(\P_mat[2][14] ) );
  GeneralPropagate_21 PM2_1_8 ( .G_ik(\G_mat[1][16] ), .P_ik(\P_mat[1][16] ), 
        .G_km1_j(\G_mat[1][15] ), .P_km1_j(\P_mat[1][15] ), .G_ij(
        \G_mat[2][16] ), .P_ij(\P_mat[2][16] ) );
  GeneralPropagate_20 PM2_1_9 ( .G_ik(\G_mat[1][18] ), .P_ik(\P_mat[1][18] ), 
        .G_km1_j(\G_mat[1][17] ), .P_km1_j(\P_mat[1][17] ), .G_ij(
        \G_mat[2][18] ), .P_ij(\P_mat[2][18] ) );
  GeneralPropagate_19 PM2_1_10 ( .G_ik(\G_mat[1][20] ), .P_ik(\P_mat[1][20] ), 
        .G_km1_j(\G_mat[1][19] ), .P_km1_j(\P_mat[1][19] ), .G_ij(
        \G_mat[2][20] ), .P_ij(\P_mat[2][20] ) );
  GeneralPropagate_18 PM2_1_11 ( .G_ik(\G_mat[1][22] ), .P_ik(\P_mat[1][22] ), 
        .G_km1_j(\G_mat[1][21] ), .P_km1_j(\P_mat[1][21] ), .G_ij(
        \G_mat[2][22] ), .P_ij(\P_mat[2][22] ) );
  GeneralPropagate_17 PM2_1_12 ( .G_ik(\G_mat[1][24] ), .P_ik(\P_mat[1][24] ), 
        .G_km1_j(\G_mat[1][23] ), .P_km1_j(\P_mat[1][23] ), .G_ij(
        \G_mat[2][24] ), .P_ij(\P_mat[2][24] ) );
  GeneralPropagate_16 PM2_1_13 ( .G_ik(\G_mat[1][26] ), .P_ik(\P_mat[1][26] ), 
        .G_km1_j(\G_mat[1][25] ), .P_km1_j(\P_mat[1][25] ), .G_ij(
        \G_mat[2][26] ), .P_ij(\P_mat[2][26] ) );
  GeneralPropagate_15 PM2_1_14 ( .G_ik(\G_mat[1][28] ), .P_ik(\P_mat[1][28] ), 
        .G_km1_j(\G_mat[1][27] ), .P_km1_j(\P_mat[1][27] ), .G_ij(
        \G_mat[2][28] ), .P_ij(\P_mat[2][28] ) );
  GeneralPropagate_14 PM2_1_15 ( .G_ik(\G_mat[1][30] ), .P_ik(\P_mat[1][30] ), 
        .G_km1_j(\G_mat[1][29] ), .P_km1_j(\P_mat[1][29] ), .G_ij(
        \G_mat[2][30] ), .P_ij(\P_mat[2][30] ) );
  GeneralPropagate_13 PM2_1_16 ( .G_ik(\G_mat[1][32] ), .P_ik(\P_mat[1][32] ), 
        .G_km1_j(\G_mat[1][31] ), .P_km1_j(\P_mat[1][31] ), .G_ij(
        \G_mat[2][32] ), .P_ij(\P_mat[2][32] ) );
  GeneralGenerate_9 PM0_2_1 ( .G_ik(\G_mat[2][4] ), .P_ik(\P_mat[2][4] ), 
        .G_km1_j(\G_mat[2][2] ), .G_ij(CarryVector[0]) );
  GeneralPropagate_12 PM2_2_2 ( .G_ik(\G_mat[2][8] ), .P_ik(\P_mat[2][8] ), 
        .G_km1_j(\G_mat[2][6] ), .P_km1_j(\P_mat[2][6] ), .G_ij(\G_mat[3][8] ), 
        .P_ij(\P_mat[3][8] ) );
  GeneralPropagate_11 PM2_2_3 ( .G_ik(\G_mat[2][12] ), .P_ik(\P_mat[2][12] ), 
        .G_km1_j(\G_mat[2][10] ), .P_km1_j(\P_mat[2][10] ), .G_ij(
        \G_mat[3][12] ), .P_ij(\P_mat[3][12] ) );
  GeneralPropagate_10 PM2_2_4 ( .G_ik(\G_mat[2][16] ), .P_ik(\P_mat[2][16] ), 
        .G_km1_j(\G_mat[2][14] ), .P_km1_j(\P_mat[2][14] ), .G_ij(
        \G_mat[3][16] ), .P_ij(\P_mat[3][16] ) );
  GeneralPropagate_9 PM2_2_5 ( .G_ik(\G_mat[2][20] ), .P_ik(\P_mat[2][20] ), 
        .G_km1_j(\G_mat[2][18] ), .P_km1_j(\P_mat[2][18] ), .G_ij(
        \G_mat[3][20] ), .P_ij(\P_mat[3][20] ) );
  GeneralPropagate_8 PM2_2_6 ( .G_ik(\G_mat[2][24] ), .P_ik(\P_mat[2][24] ), 
        .G_km1_j(\G_mat[2][22] ), .P_km1_j(\P_mat[2][22] ), .G_ij(
        \G_mat[3][24] ), .P_ij(\P_mat[3][24] ) );
  GeneralPropagate_7 PM2_2_7 ( .G_ik(\G_mat[2][28] ), .P_ik(\P_mat[2][28] ), 
        .G_km1_j(\G_mat[2][26] ), .P_km1_j(\P_mat[2][26] ), .G_ij(
        \G_mat[3][28] ), .P_ij(\P_mat[3][28] ) );
  GeneralPropagate_6 PM2_2_8 ( .G_ik(\G_mat[2][32] ), .P_ik(\P_mat[2][32] ), 
        .G_km1_j(\G_mat[2][30] ), .P_km1_j(\P_mat[2][30] ), .G_ij(
        \G_mat[3][32] ), .P_ij(\P_mat[3][32] ) );
  GeneralGenerate_8 PM0_3_1 ( .G_ik(\G_mat[3][8] ), .P_ik(\P_mat[3][8] ), 
        .G_km1_j(CarryVector[0]), .G_ij(CarryVector[1]) );
  GeneralPropagate_5 PM2_3_2 ( .G_ik(\G_mat[3][16] ), .P_ik(\P_mat[3][16] ), 
        .G_km1_j(\G_mat[3][12] ), .P_km1_j(\P_mat[3][12] ), .G_ij(
        \G_mat[4][16] ), .P_ij(\P_mat[4][16] ) );
  GeneralPropagate_4 PM2_3_3 ( .G_ik(\G_mat[3][24] ), .P_ik(\P_mat[3][24] ), 
        .G_km1_j(\G_mat[3][20] ), .P_km1_j(\P_mat[3][20] ), .G_ij(
        \G_mat[4][24] ), .P_ij(\P_mat[4][24] ) );
  GeneralPropagate_3 PM2_3_4 ( .G_ik(\G_mat[3][32] ), .P_ik(\P_mat[3][32] ), 
        .G_km1_j(\G_mat[3][28] ), .P_km1_j(\P_mat[3][28] ), .G_ij(
        \G_mat[4][32] ), .P_ij(\P_mat[4][32] ) );
  GeneralGenerate_7 PM3_4_1_1 ( .G_ik(\G_mat[4][16] ), .P_ik(\P_mat[4][16] ), 
        .G_km1_j(CarryVector[1]), .G_ij(CarryVector[3]) );
  GeneralGenerate_6 PM4_4_1_1 ( .G_ik(\G_mat[3][12] ), .P_ik(\P_mat[3][12] ), 
        .G_km1_j(CarryVector[1]), .G_ij(CarryVector[2]) );
  GeneralPropagate_2 PM7_4_2_1 ( .G_ik(\G_mat[4][32] ), .P_ik(\P_mat[4][32] ), 
        .G_km1_j(\G_mat[4][24] ), .P_km1_j(\P_mat[4][24] ), .G_ij(
        \G_mat[5][32] ), .P_ij(\P_mat[5][32] ) );
  GeneralPropagate_1 PM5_4_2_1 ( .G_ik(\G_mat[3][28] ), .P_ik(\P_mat[3][28] ), 
        .G_km1_j(\G_mat[4][24] ), .P_km1_j(\P_mat[4][24] ), .G_ij(
        \G_mat[5][28] ), .P_ij(\P_mat[5][28] ) );
  GeneralGenerate_5 PM9_5_1 ( .G_ik(\G_mat[5][32] ), .P_ik(\P_mat[5][32] ), 
        .G_km1_j(CarryVector[3]), .G_ij(CarryVector[7]) );
  GeneralGenerate_4 PM9_5_2 ( .G_ik(\G_mat[5][28] ), .P_ik(\P_mat[5][28] ), 
        .G_km1_j(CarryVector[3]), .G_ij(CarryVector[6]) );
  GeneralGenerate_3 PM14_5_1_1 ( .G_ik(\G_mat[4][24] ), .P_ik(\P_mat[4][24] ), 
        .G_km1_j(CarryVector[3]), .G_ij(CarryVector[5]) );
  GeneralGenerate_2 PM13_5_2 ( .G_ik(\G_mat[3][20] ), .P_ik(\P_mat[3][20] ), 
        .G_km1_j(CarryVector[3]), .G_ij(CarryVector[4]) );
endmodule


module Mux_NBit_2x1_NBIT_IN3 ( port0, port1, sel, portY );
  input [2:0] port0;
  input [2:0] port1;
  output [2:0] portY;
  input sel;
  wire   N2, N4, n5, n7, n8, n2;
  assign portY[0] = N2;
  assign portY[2] = N4;

  INV_X1 U1 ( .A(n8), .ZN(N2) );
  AOI22_X1 U2 ( .A1(port0[0]), .A2(n2), .B1(port1[0]), .B2(sel), .ZN(n8) );
  INV_X1 U3 ( .A(n5), .ZN(portY[1]) );
  AOI22_X1 U4 ( .A1(port0[1]), .A2(n2), .B1(sel), .B2(port1[1]), .ZN(n5) );
  INV_X1 U5 ( .A(n7), .ZN(N4) );
  AOI22_X1 U6 ( .A1(port0[2]), .A2(n2), .B1(port1[2]), .B2(sel), .ZN(n7) );
  INV_X1 U7 ( .A(sel), .ZN(n2) );
endmodule


module Mux_NBit_2x1_NBIT_IN40_1 ( port0, port1, sel, portY );
  input [39:0] port0;
  input [39:0] port1;
  output [39:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, n42, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n57, n58, n59, n60, n61,
         n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;
  assign portY[32] = N34;
  assign portY[33] = N35;
  assign portY[34] = N36;
  assign portY[35] = N37;
  assign portY[36] = N38;
  assign portY[37] = N39;
  assign portY[38] = N40;
  assign portY[39] = N41;

  INV_X2 U41 ( .A(n63), .ZN(N28) );
  MUX2_X2 U1 ( .A(port0[33]), .B(port1[33]), .S(sel), .Z(N35) );
  MUX2_X2 U2 ( .A(port0[32]), .B(port1[32]), .S(sel), .Z(N34) );
  INV_X1 U3 ( .A(n62), .ZN(N29) );
  INV_X1 U4 ( .A(n58), .ZN(N32) );
  INV_X1 U5 ( .A(n66), .ZN(N25) );
  INV_X1 U6 ( .A(n65), .ZN(N26) );
  INV_X1 U7 ( .A(n59), .ZN(N31) );
  INV_X1 U8 ( .A(n60), .ZN(N30) );
  BUF_X1 U9 ( .A(n8), .Z(n23) );
  CLKBUF_X1 U10 ( .A(n6), .Z(n17) );
  CLKBUF_X1 U11 ( .A(n9), .Z(n7) );
  INV_X1 U12 ( .A(n23), .ZN(n12) );
  INV_X1 U13 ( .A(n23), .ZN(n11) );
  BUF_X1 U14 ( .A(n7), .Z(n20) );
  BUF_X1 U15 ( .A(n7), .Z(n19) );
  BUF_X1 U16 ( .A(n6), .Z(n18) );
  BUF_X1 U17 ( .A(n5), .Z(n14) );
  BUF_X1 U18 ( .A(n6), .Z(n16) );
  BUF_X1 U19 ( .A(n5), .Z(n15) );
  BUF_X1 U20 ( .A(n7), .Z(n21) );
  CLKBUF_X1 U21 ( .A(n8), .Z(n22) );
  CLKBUF_X1 U22 ( .A(n5), .Z(n13) );
  BUF_X1 U23 ( .A(n10), .Z(n6) );
  BUF_X1 U24 ( .A(n10), .Z(n5) );
  BUF_X1 U25 ( .A(n9), .Z(n8) );
  CLKBUF_X1 U26 ( .A(sel), .Z(n9) );
  CLKBUF_X1 U27 ( .A(sel), .Z(n10) );
  AOI22_X1 U28 ( .A1(port0[29]), .A2(n12), .B1(port1[29]), .B2(n16), .ZN(n59)
         );
  AOI22_X1 U29 ( .A1(port0[28]), .A2(n12), .B1(port1[28]), .B2(n16), .ZN(n60)
         );
  AOI22_X1 U30 ( .A1(port0[37]), .A2(n11), .B1(port1[37]), .B2(n14), .ZN(n51)
         );
  AOI22_X1 U31 ( .A1(port0[36]), .A2(n12), .B1(port1[36]), .B2(n15), .ZN(n52)
         );
  INV_X1 U32 ( .A(n48), .ZN(N41) );
  AOI22_X1 U33 ( .A1(port0[39]), .A2(n12), .B1(port1[39]), .B2(n14), .ZN(n48)
         );
  INV_X1 U34 ( .A(n64), .ZN(N27) );
  AOI22_X1 U35 ( .A1(port0[25]), .A2(n12), .B1(port1[25]), .B2(n17), .ZN(n64)
         );
  AOI22_X1 U36 ( .A1(port0[27]), .A2(n12), .B1(port1[27]), .B2(n17), .ZN(n62)
         );
  AOI22_X1 U37 ( .A1(port0[26]), .A2(n12), .B1(port1[26]), .B2(n17), .ZN(n63)
         );
  INV_X1 U38 ( .A(n76), .ZN(N16) );
  AOI22_X1 U39 ( .A1(port0[14]), .A2(n11), .B1(port1[14]), .B2(n21), .ZN(n76)
         );
  AOI22_X1 U40 ( .A1(port0[24]), .A2(n12), .B1(port1[24]), .B2(n18), .ZN(n65)
         );
  AOI22_X1 U42 ( .A1(port0[23]), .A2(n12), .B1(port1[23]), .B2(n18), .ZN(n66)
         );
  INV_X1 U43 ( .A(n67), .ZN(N24) );
  AOI22_X1 U44 ( .A1(port0[22]), .A2(n12), .B1(port1[22]), .B2(n18), .ZN(n67)
         );
  INV_X1 U45 ( .A(n70), .ZN(N21) );
  AOI22_X1 U46 ( .A1(port0[19]), .A2(n12), .B1(port1[19]), .B2(n19), .ZN(n70)
         );
  INV_X1 U47 ( .A(n69), .ZN(N22) );
  AOI22_X1 U48 ( .A1(port0[20]), .A2(n12), .B1(port1[20]), .B2(n19), .ZN(n69)
         );
  INV_X1 U49 ( .A(n68), .ZN(N23) );
  AOI22_X1 U50 ( .A1(port0[21]), .A2(n12), .B1(port1[21]), .B2(n19), .ZN(n68)
         );
  INV_X1 U51 ( .A(n73), .ZN(N19) );
  AOI22_X1 U52 ( .A1(port0[17]), .A2(n11), .B1(port1[17]), .B2(n20), .ZN(n73)
         );
  INV_X1 U53 ( .A(n71), .ZN(N20) );
  AOI22_X1 U54 ( .A1(port0[18]), .A2(n11), .B1(port1[18]), .B2(n19), .ZN(n71)
         );
  INV_X1 U55 ( .A(n75), .ZN(N17) );
  AOI22_X1 U56 ( .A1(port0[15]), .A2(n11), .B1(port1[15]), .B2(n20), .ZN(n75)
         );
  INV_X1 U57 ( .A(n77), .ZN(N15) );
  AOI22_X1 U58 ( .A1(port0[13]), .A2(n11), .B1(port1[13]), .B2(n21), .ZN(n77)
         );
  INV_X1 U59 ( .A(n80), .ZN(N12) );
  AOI22_X1 U60 ( .A1(port0[10]), .A2(n11), .B1(port1[10]), .B2(n22), .ZN(n80)
         );
  INV_X1 U61 ( .A(n78), .ZN(N14) );
  AOI22_X1 U62 ( .A1(port0[12]), .A2(n11), .B1(port1[12]), .B2(n21), .ZN(n78)
         );
  INV_X1 U63 ( .A(n79), .ZN(N13) );
  AOI22_X1 U64 ( .A1(port0[11]), .A2(n11), .B1(port1[11]), .B2(n21), .ZN(n79)
         );
  INV_X1 U65 ( .A(n74), .ZN(N18) );
  AOI22_X1 U66 ( .A1(port0[16]), .A2(n11), .B1(port1[16]), .B2(n20), .ZN(n74)
         );
  INV_X1 U67 ( .A(n82), .ZN(N10) );
  AOI22_X1 U68 ( .A1(port0[8]), .A2(n11), .B1(port1[8]), .B2(n22), .ZN(n82) );
  INV_X1 U69 ( .A(n81), .ZN(N11) );
  AOI22_X1 U70 ( .A1(port0[9]), .A2(n11), .B1(port1[9]), .B2(n22), .ZN(n81) );
  INV_X1 U71 ( .A(n42), .ZN(N9) );
  AOI22_X1 U72 ( .A1(port0[7]), .A2(n11), .B1(n22), .B2(port1[7]), .ZN(n42) );
  INV_X1 U73 ( .A(n44), .ZN(N8) );
  AOI22_X1 U74 ( .A1(port0[6]), .A2(n11), .B1(port1[6]), .B2(n13), .ZN(n44) );
  INV_X1 U75 ( .A(n61), .ZN(N3) );
  AOI22_X1 U76 ( .A1(port0[1]), .A2(n12), .B1(port1[1]), .B2(n17), .ZN(n61) );
  INV_X1 U77 ( .A(n45), .ZN(N7) );
  AOI22_X1 U78 ( .A1(port0[5]), .A2(n11), .B1(port1[5]), .B2(n13), .ZN(n45) );
  INV_X1 U79 ( .A(n46), .ZN(N6) );
  AOI22_X1 U80 ( .A1(port0[4]), .A2(n11), .B1(port1[4]), .B2(n13), .ZN(n46) );
  INV_X1 U81 ( .A(n47), .ZN(N5) );
  AOI22_X1 U82 ( .A1(port0[3]), .A2(n11), .B1(port1[3]), .B2(n13), .ZN(n47) );
  INV_X1 U83 ( .A(n50), .ZN(N4) );
  AOI22_X1 U84 ( .A1(port0[2]), .A2(n12), .B1(port1[2]), .B2(n14), .ZN(n50) );
  INV_X1 U85 ( .A(n72), .ZN(N2) );
  AOI22_X1 U86 ( .A1(port0[0]), .A2(n11), .B1(port1[0]), .B2(n20), .ZN(n72) );
  AOI22_X1 U87 ( .A1(port0[30]), .A2(n11), .B1(port1[30]), .B2(n16), .ZN(n58)
         );
  INV_X1 U88 ( .A(n49), .ZN(N40) );
  AOI22_X1 U89 ( .A1(port0[35]), .A2(n12), .B1(port1[35]), .B2(n18), .ZN(n53)
         );
  AOI22_X1 U90 ( .A1(port0[38]), .A2(n12), .B1(port1[38]), .B2(n14), .ZN(n49)
         );
  INV_X1 U91 ( .A(n51), .ZN(N39) );
  INV_X1 U92 ( .A(n57), .ZN(N33) );
  INV_X1 U93 ( .A(n53), .ZN(N37) );
  AOI22_X1 U94 ( .A1(port0[31]), .A2(n11), .B1(port1[31]), .B2(n16), .ZN(n57)
         );
  INV_X1 U95 ( .A(n52), .ZN(N38) );
  INV_X1 U96 ( .A(n54), .ZN(N36) );
  AOI22_X1 U97 ( .A1(port0[34]), .A2(n12), .B1(port1[34]), .B2(n15), .ZN(n54)
         );
endmodule


module Mux_NBit_2x1_NBIT_IN40_0 ( port0, port1, sel, portY );
  input [39:0] port0;
  input [39:0] port1;
  output [39:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, n42, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73,
         n74, n75, n76, n77, n78, n79, n80, n81, n82, n1, n2, n3, n4, n5, n6,
         n7, n8, n9, n10, n11, n12, n13;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;
  assign portY[32] = N34;
  assign portY[33] = N35;
  assign portY[34] = N36;
  assign portY[35] = N37;
  assign portY[36] = N38;
  assign portY[37] = N39;
  assign portY[38] = N40;
  assign portY[39] = N41;

  CLKBUF_X1 U1 ( .A(sel), .Z(n1) );
  BUF_X2 U2 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U3 ( .A(n2), .Z(n11) );
  INV_X1 U4 ( .A(n3), .ZN(n5) );
  INV_X1 U5 ( .A(n3), .ZN(n4) );
  BUF_X1 U6 ( .A(n2), .Z(n12) );
  BUF_X1 U7 ( .A(n2), .Z(n10) );
  BUF_X1 U8 ( .A(n1), .Z(n9) );
  BUF_X1 U9 ( .A(n1), .Z(n8) );
  AOI22_X1 U10 ( .A1(port0[23]), .A2(n6), .B1(port1[23]), .B2(n12), .ZN(n66)
         );
  AOI22_X1 U11 ( .A1(port0[16]), .A2(n6), .B1(port1[16]), .B2(n13), .ZN(n74)
         );
  AOI22_X1 U12 ( .A1(port0[22]), .A2(n7), .B1(port1[22]), .B2(n12), .ZN(n67)
         );
  AOI22_X1 U13 ( .A1(port0[21]), .A2(n4), .B1(port1[21]), .B2(n13), .ZN(n68)
         );
  AOI22_X1 U14 ( .A1(port0[20]), .A2(n6), .B1(port1[20]), .B2(n13), .ZN(n69)
         );
  AOI22_X1 U15 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n71)
         );
  AOI22_X1 U16 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n13), .ZN(n73)
         );
  AOI22_X1 U17 ( .A1(port0[19]), .A2(n6), .B1(port1[19]), .B2(n13), .ZN(n70)
         );
  CLKBUF_X1 U18 ( .A(n3), .Z(n13) );
  INV_X1 U19 ( .A(n55), .ZN(N35) );
  AOI22_X1 U20 ( .A1(port0[27]), .A2(n6), .B1(port1[27]), .B2(n11), .ZN(n62)
         );
  AOI22_X1 U21 ( .A1(port0[26]), .A2(n7), .B1(port1[26]), .B2(n11), .ZN(n63)
         );
  AOI22_X1 U22 ( .A1(port0[25]), .A2(n4), .B1(port1[25]), .B2(n11), .ZN(n64)
         );
  INV_X1 U23 ( .A(n60), .ZN(N30) );
  INV_X1 U24 ( .A(n62), .ZN(N29) );
  INV_X1 U25 ( .A(n64), .ZN(N27) );
  INV_X1 U26 ( .A(n59), .ZN(N31) );
  INV_X1 U27 ( .A(n49), .ZN(N40) );
  BUF_X1 U28 ( .A(sel), .Z(n2) );
  INV_X1 U29 ( .A(n51), .ZN(N39) );
  INV_X1 U30 ( .A(n53), .ZN(N37) );
  INV_X1 U31 ( .A(n48), .ZN(N41) );
  AOI22_X1 U32 ( .A1(port0[24]), .A2(n6), .B1(port1[24]), .B2(n12), .ZN(n65)
         );
  INV_X1 U33 ( .A(n65), .ZN(N26) );
  AOI22_X1 U34 ( .A1(port0[29]), .A2(n7), .B1(port1[29]), .B2(n10), .ZN(n59)
         );
  AOI22_X1 U35 ( .A1(port0[28]), .A2(n6), .B1(port1[28]), .B2(n10), .ZN(n60)
         );
  INV_X1 U36 ( .A(n63), .ZN(N28) );
  AOI22_X1 U37 ( .A1(port0[15]), .A2(n6), .B1(port1[15]), .B2(n13), .ZN(n75)
         );
  AOI22_X1 U38 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n13), .ZN(n76)
         );
  AOI22_X1 U39 ( .A1(port0[9]), .A2(n6), .B1(port1[9]), .B2(n13), .ZN(n81) );
  AOI22_X1 U40 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n13), .ZN(n80)
         );
  AOI22_X1 U41 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n13), .ZN(n77)
         );
  AOI22_X1 U42 ( .A1(port0[12]), .A2(n6), .B1(port1[12]), .B2(n13), .ZN(n78)
         );
  AOI22_X1 U43 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n13), .ZN(n79)
         );
  INV_X1 U44 ( .A(n67), .ZN(N24) );
  INV_X1 U45 ( .A(n69), .ZN(N22) );
  INV_X1 U46 ( .A(n68), .ZN(N23) );
  INV_X1 U47 ( .A(n74), .ZN(N18) );
  INV_X1 U48 ( .A(n71), .ZN(N20) );
  INV_X1 U49 ( .A(n73), .ZN(N19) );
  INV_X1 U50 ( .A(n75), .ZN(N17) );
  INV_X1 U51 ( .A(n76), .ZN(N16) );
  INV_X1 U52 ( .A(n80), .ZN(N12) );
  INV_X1 U53 ( .A(n77), .ZN(N15) );
  INV_X1 U54 ( .A(n78), .ZN(N14) );
  INV_X1 U55 ( .A(n79), .ZN(N13) );
  INV_X1 U56 ( .A(n66), .ZN(N25) );
  INV_X1 U57 ( .A(n70), .ZN(N21) );
  INV_X1 U58 ( .A(n81), .ZN(N11) );
  AOI22_X1 U59 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n82) );
  INV_X1 U60 ( .A(n72), .ZN(N2) );
  INV_X1 U61 ( .A(n82), .ZN(N10) );
  INV_X1 U62 ( .A(n47), .ZN(N5) );
  INV_X1 U63 ( .A(n50), .ZN(N4) );
  INV_X1 U64 ( .A(n61), .ZN(N3) );
  INV_X1 U65 ( .A(n42), .ZN(N9) );
  INV_X1 U66 ( .A(n44), .ZN(N8) );
  INV_X1 U67 ( .A(n45), .ZN(N7) );
  INV_X1 U68 ( .A(n46), .ZN(N6) );
  AOI22_X1 U69 ( .A1(port0[1]), .A2(n4), .B1(port1[1]), .B2(n11), .ZN(n61) );
  AOI22_X1 U70 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n13), .ZN(n72) );
  AOI22_X1 U71 ( .A1(port0[7]), .A2(n7), .B1(n13), .B2(port1[7]), .ZN(n42) );
  AOI22_X1 U72 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n8), .ZN(n44) );
  AOI22_X1 U73 ( .A1(port0[5]), .A2(n6), .B1(port1[5]), .B2(n13), .ZN(n45) );
  AOI22_X1 U74 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n8), .ZN(n46) );
  AOI22_X1 U75 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n8), .ZN(n50) );
  AOI22_X1 U76 ( .A1(port0[3]), .A2(n7), .B1(port1[3]), .B2(n13), .ZN(n47) );
  AOI22_X1 U77 ( .A1(port0[39]), .A2(n4), .B1(port1[39]), .B2(n8), .ZN(n48) );
  AOI22_X1 U78 ( .A1(port0[38]), .A2(n4), .B1(port1[38]), .B2(n3), .ZN(n49) );
  AOI22_X1 U79 ( .A1(port0[37]), .A2(n7), .B1(port1[37]), .B2(n8), .ZN(n51) );
  AOI22_X1 U80 ( .A1(port0[36]), .A2(n6), .B1(port1[36]), .B2(n8), .ZN(n52) );
  AOI22_X1 U81 ( .A1(port0[34]), .A2(n5), .B1(port1[34]), .B2(n9), .ZN(n54) );
  AOI22_X1 U82 ( .A1(port0[35]), .A2(n5), .B1(port1[35]), .B2(n12), .ZN(n53)
         );
  AOI22_X1 U83 ( .A1(port0[32]), .A2(n5), .B1(port1[32]), .B2(n9), .ZN(n56) );
  AOI22_X1 U84 ( .A1(port0[31]), .A2(n5), .B1(port1[31]), .B2(n10), .ZN(n57)
         );
  INV_X1 U85 ( .A(n52), .ZN(N38) );
  INV_X1 U86 ( .A(n58), .ZN(N32) );
  AOI22_X1 U87 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n10), .ZN(n58)
         );
  INV_X1 U88 ( .A(n54), .ZN(N36) );
  INV_X1 U89 ( .A(n56), .ZN(N34) );
  INV_X1 U90 ( .A(n57), .ZN(N33) );
  AOI22_X1 U91 ( .A1(port0[33]), .A2(n5), .B1(port1[33]), .B2(n9), .ZN(n55) );
  INV_X2 U92 ( .A(n3), .ZN(n6) );
  INV_X1 U93 ( .A(n3), .ZN(n7) );
endmodule


module Mux_NBit_2x1_NBIT_IN8_0 ( port0, port1, sel, portY );
  input [7:0] port0;
  input [7:0] port1;
  output [7:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, n11, n12, n13, n14, n16;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;

  MUX2_X2 U1 ( .A(port1[1]), .B(port0[1]), .S(n11), .Z(N3) );
  MUX2_X1 U2 ( .A(port0[7]), .B(port1[7]), .S(sel), .Z(N9) );
  MUX2_X1 U3 ( .A(port0[3]), .B(port1[3]), .S(sel), .Z(N5) );
  MUX2_X1 U4 ( .A(port0[0]), .B(port1[0]), .S(sel), .Z(N2) );
  INV_X1 U5 ( .A(sel), .ZN(n11) );
  INV_X1 U6 ( .A(n13), .ZN(N7) );
  INV_X1 U7 ( .A(n14), .ZN(N6) );
  INV_X1 U8 ( .A(n12), .ZN(N8) );
  INV_X1 U9 ( .A(n16), .ZN(N4) );
  AOI22_X1 U10 ( .A1(port0[5]), .A2(n11), .B1(port1[5]), .B2(sel), .ZN(n13) );
  AOI22_X1 U11 ( .A1(port0[6]), .A2(n11), .B1(port1[6]), .B2(sel), .ZN(n12) );
  AOI22_X1 U12 ( .A1(port0[4]), .A2(n11), .B1(port1[4]), .B2(sel), .ZN(n14) );
  AOI22_X1 U13 ( .A1(port0[2]), .A2(n11), .B1(port1[2]), .B2(sel), .ZN(n16) );
endmodule


module PG_cell_0 ( A, B, p, g );
  input A, B;
  output p, g;


  XOR2_X1 U2 ( .A(B), .B(A), .Z(p) );
  AND2_X1 U1 ( .A1(B), .A2(A), .ZN(g) );
endmodule


module GeneralGenerate_0 ( G_ik, P_ik, G_km1_j, G_ij );
  input G_ik, P_ik, G_km1_j;
  output G_ij;
  wire   n2;

  INV_X1 U1 ( .A(n2), .ZN(G_ij) );
  AOI21_X1 U2 ( .B1(P_ik), .B2(G_km1_j), .A(G_ik), .ZN(n2) );
endmodule


module t_ff_rst1_32 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFS_X1 data_reg ( .D(n3), .CK(TFF_clk), .SN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_64 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n3, n4;

  DFFR_X1 data_reg ( .D(n3), .CK(TFF_clk), .RN(n4), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n3) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n4) );
endmodule


module t_ff_rst0_0 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n1, n2;

  DFFR_X1 data_reg ( .D(n2), .CK(TFF_clk), .RN(n1), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n2) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n1) );
endmodule


module t_ff_rst1_0 ( TFF_clk, TFF_rst, TFF_t, TFF_q, TFF_nq );
  input TFF_clk, TFF_rst, TFF_t;
  output TFF_q, TFF_nq;
  wire   n1, n2;

  DFFS_X1 data_reg ( .D(n2), .CK(TFF_clk), .SN(n1), .Q(TFF_q), .QN(TFF_nq) );
  XOR2_X1 U3 ( .A(TFF_t), .B(TFF_q), .Z(n2) );
  INV_X1 U2 ( .A(TFF_rst), .ZN(n1) );
endmodule


module Multiplier_NBIT_DATA32_DW02_mult_1 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   \ab[31][31] , \ab[31][30] , \ab[31][29] , \ab[31][28] , \ab[31][27] ,
         \ab[31][26] , \ab[31][25] , \ab[31][24] , \ab[31][23] , \ab[31][22] ,
         \ab[31][21] , \ab[31][20] , \ab[31][19] , \ab[31][18] , \ab[31][17] ,
         \ab[31][16] , \ab[31][15] , \ab[31][14] , \ab[31][13] , \ab[31][12] ,
         \ab[31][11] , \ab[31][10] , \ab[31][9] , \ab[31][8] , \ab[31][7] ,
         \ab[31][6] , \ab[31][5] , \ab[31][4] , \ab[31][3] , \ab[31][2] ,
         \ab[31][1] , \ab[31][0] , \ab[30][31] , \ab[30][30] , \ab[30][29] ,
         \ab[30][28] , \ab[30][27] , \ab[30][26] , \ab[30][25] , \ab[30][24] ,
         \ab[30][23] , \ab[30][22] , \ab[30][21] , \ab[30][20] , \ab[30][19] ,
         \ab[30][18] , \ab[30][17] , \ab[30][16] , \ab[30][15] , \ab[30][14] ,
         \ab[30][13] , \ab[30][12] , \ab[30][11] , \ab[30][10] , \ab[30][9] ,
         \ab[30][8] , \ab[30][7] , \ab[30][6] , \ab[30][5] , \ab[30][4] ,
         \ab[30][3] , \ab[30][2] , \ab[30][1] , \ab[30][0] , \ab[29][31] ,
         \ab[29][30] , \ab[29][29] , \ab[29][28] , \ab[29][27] , \ab[29][26] ,
         \ab[29][25] , \ab[29][24] , \ab[29][23] , \ab[29][22] , \ab[29][21] ,
         \ab[29][20] , \ab[29][19] , \ab[29][18] , \ab[29][17] , \ab[29][16] ,
         \ab[29][15] , \ab[29][14] , \ab[29][13] , \ab[29][12] , \ab[29][11] ,
         \ab[29][10] , \ab[29][9] , \ab[29][8] , \ab[29][7] , \ab[29][6] ,
         \ab[29][5] , \ab[29][4] , \ab[29][3] , \ab[29][2] , \ab[29][1] ,
         \ab[29][0] , \ab[28][31] , \ab[28][30] , \ab[28][29] , \ab[28][28] ,
         \ab[28][27] , \ab[28][26] , \ab[28][25] , \ab[28][24] , \ab[28][23] ,
         \ab[28][22] , \ab[28][21] , \ab[28][20] , \ab[28][19] , \ab[28][18] ,
         \ab[28][17] , \ab[28][16] , \ab[28][15] , \ab[28][14] , \ab[28][13] ,
         \ab[28][12] , \ab[28][11] , \ab[28][10] , \ab[28][9] , \ab[28][8] ,
         \ab[28][7] , \ab[28][6] , \ab[28][5] , \ab[28][4] , \ab[28][3] ,
         \ab[28][2] , \ab[28][1] , \ab[28][0] , \ab[27][31] , \ab[27][30] ,
         \ab[27][29] , \ab[27][28] , \ab[27][27] , \ab[27][26] , \ab[27][25] ,
         \ab[27][24] , \ab[27][23] , \ab[27][22] , \ab[27][21] , \ab[27][20] ,
         \ab[27][19] , \ab[27][18] , \ab[27][17] , \ab[27][16] , \ab[27][15] ,
         \ab[27][14] , \ab[27][13] , \ab[27][12] , \ab[27][11] , \ab[27][10] ,
         \ab[27][9] , \ab[27][8] , \ab[27][7] , \ab[27][6] , \ab[27][5] ,
         \ab[27][4] , \ab[27][3] , \ab[27][2] , \ab[27][1] , \ab[27][0] ,
         \ab[26][31] , \ab[26][30] , \ab[26][29] , \ab[26][28] , \ab[26][27] ,
         \ab[26][26] , \ab[26][25] , \ab[26][24] , \ab[26][23] , \ab[26][22] ,
         \ab[26][21] , \ab[26][20] , \ab[26][19] , \ab[26][18] , \ab[26][17] ,
         \ab[26][16] , \ab[26][15] , \ab[26][14] , \ab[26][13] , \ab[26][12] ,
         \ab[26][11] , \ab[26][10] , \ab[26][9] , \ab[26][8] , \ab[26][7] ,
         \ab[26][6] , \ab[26][5] , \ab[26][4] , \ab[26][3] , \ab[26][2] ,
         \ab[26][1] , \ab[26][0] , \ab[25][31] , \ab[25][30] , \ab[25][29] ,
         \ab[25][28] , \ab[25][27] , \ab[25][26] , \ab[25][25] , \ab[25][24] ,
         \ab[25][23] , \ab[25][22] , \ab[25][21] , \ab[25][20] , \ab[25][19] ,
         \ab[25][18] , \ab[25][17] , \ab[25][16] , \ab[25][15] , \ab[25][14] ,
         \ab[25][13] , \ab[25][12] , \ab[25][11] , \ab[25][10] , \ab[25][9] ,
         \ab[25][8] , \ab[25][7] , \ab[25][6] , \ab[25][5] , \ab[25][4] ,
         \ab[25][3] , \ab[25][2] , \ab[25][1] , \ab[25][0] , \ab[24][31] ,
         \ab[24][30] , \ab[24][29] , \ab[24][28] , \ab[24][27] , \ab[24][26] ,
         \ab[24][25] , \ab[24][24] , \ab[24][23] , \ab[24][22] , \ab[24][21] ,
         \ab[24][20] , \ab[24][19] , \ab[24][18] , \ab[24][17] , \ab[24][16] ,
         \ab[24][15] , \ab[24][14] , \ab[24][13] , \ab[24][12] , \ab[24][11] ,
         \ab[24][10] , \ab[24][9] , \ab[24][8] , \ab[24][7] , \ab[24][6] ,
         \ab[24][5] , \ab[24][4] , \ab[24][3] , \ab[24][2] , \ab[24][1] ,
         \ab[24][0] , \ab[23][31] , \ab[23][30] , \ab[23][29] , \ab[23][28] ,
         \ab[23][27] , \ab[23][26] , \ab[23][25] , \ab[23][24] , \ab[23][23] ,
         \ab[23][22] , \ab[23][21] , \ab[23][20] , \ab[23][19] , \ab[23][18] ,
         \ab[23][17] , \ab[23][16] , \ab[23][15] , \ab[23][14] , \ab[23][13] ,
         \ab[23][12] , \ab[23][11] , \ab[23][10] , \ab[23][9] , \ab[23][8] ,
         \ab[23][7] , \ab[23][6] , \ab[23][5] , \ab[23][4] , \ab[23][3] ,
         \ab[23][2] , \ab[23][1] , \ab[23][0] , \ab[22][31] , \ab[22][30] ,
         \ab[22][29] , \ab[22][28] , \ab[22][27] , \ab[22][26] , \ab[22][25] ,
         \ab[22][24] , \ab[22][23] , \ab[22][22] , \ab[22][21] , \ab[22][20] ,
         \ab[22][19] , \ab[22][18] , \ab[22][17] , \ab[22][16] , \ab[22][15] ,
         \ab[22][14] , \ab[22][13] , \ab[22][12] , \ab[22][11] , \ab[22][10] ,
         \ab[22][9] , \ab[22][8] , \ab[22][7] , \ab[22][6] , \ab[22][5] ,
         \ab[22][4] , \ab[22][3] , \ab[22][2] , \ab[22][1] , \ab[22][0] ,
         \ab[21][31] , \ab[21][30] , \ab[21][29] , \ab[21][28] , \ab[21][27] ,
         \ab[21][26] , \ab[21][25] , \ab[21][24] , \ab[21][23] , \ab[21][22] ,
         \ab[21][21] , \ab[21][20] , \ab[21][19] , \ab[21][18] , \ab[21][17] ,
         \ab[21][16] , \ab[21][15] , \ab[21][14] , \ab[21][13] , \ab[21][12] ,
         \ab[21][11] , \ab[21][10] , \ab[21][9] , \ab[21][8] , \ab[21][7] ,
         \ab[21][6] , \ab[21][5] , \ab[21][4] , \ab[21][3] , \ab[21][2] ,
         \ab[21][1] , \ab[21][0] , \ab[20][31] , \ab[20][30] , \ab[20][29] ,
         \ab[20][28] , \ab[20][27] , \ab[20][26] , \ab[20][25] , \ab[20][24] ,
         \ab[20][23] , \ab[20][22] , \ab[20][21] , \ab[20][20] , \ab[20][19] ,
         \ab[20][18] , \ab[20][17] , \ab[20][16] , \ab[20][15] , \ab[20][14] ,
         \ab[20][13] , \ab[20][12] , \ab[20][11] , \ab[20][10] , \ab[20][9] ,
         \ab[20][8] , \ab[20][7] , \ab[20][6] , \ab[20][5] , \ab[20][4] ,
         \ab[20][3] , \ab[20][2] , \ab[20][1] , \ab[20][0] , \ab[19][31] ,
         \ab[19][30] , \ab[19][29] , \ab[19][28] , \ab[19][27] , \ab[19][26] ,
         \ab[19][25] , \ab[19][24] , \ab[19][23] , \ab[19][22] , \ab[19][21] ,
         \ab[19][20] , \ab[19][19] , \ab[19][18] , \ab[19][17] , \ab[19][16] ,
         \ab[19][15] , \ab[19][14] , \ab[19][13] , \ab[19][12] , \ab[19][11] ,
         \ab[19][10] , \ab[19][9] , \ab[19][8] , \ab[19][7] , \ab[19][6] ,
         \ab[19][5] , \ab[19][4] , \ab[19][3] , \ab[19][2] , \ab[19][1] ,
         \ab[19][0] , \ab[18][31] , \ab[18][30] , \ab[18][29] , \ab[18][28] ,
         \ab[18][27] , \ab[18][26] , \ab[18][25] , \ab[18][24] , \ab[18][23] ,
         \ab[18][22] , \ab[18][21] , \ab[18][20] , \ab[18][19] , \ab[18][18] ,
         \ab[18][17] , \ab[18][16] , \ab[18][15] , \ab[18][14] , \ab[18][13] ,
         \ab[18][12] , \ab[18][11] , \ab[18][10] , \ab[18][9] , \ab[18][8] ,
         \ab[18][7] , \ab[18][6] , \ab[18][5] , \ab[18][4] , \ab[18][3] ,
         \ab[18][2] , \ab[18][1] , \ab[18][0] , \ab[17][31] , \ab[17][30] ,
         \ab[17][29] , \ab[17][28] , \ab[17][27] , \ab[17][26] , \ab[17][25] ,
         \ab[17][24] , \ab[17][23] , \ab[17][22] , \ab[17][21] , \ab[17][20] ,
         \ab[17][19] , \ab[17][18] , \ab[17][17] , \ab[17][16] , \ab[17][15] ,
         \ab[17][14] , \ab[17][13] , \ab[17][12] , \ab[17][11] , \ab[17][10] ,
         \ab[17][9] , \ab[17][8] , \ab[17][7] , \ab[17][6] , \ab[17][5] ,
         \ab[17][4] , \ab[17][3] , \ab[17][2] , \ab[17][1] , \ab[17][0] ,
         \ab[16][31] , \ab[16][30] , \ab[16][29] , \ab[16][28] , \ab[16][27] ,
         \ab[16][26] , \ab[16][25] , \ab[16][24] , \ab[16][23] , \ab[16][22] ,
         \ab[16][21] , \ab[16][20] , \ab[16][19] , \ab[16][18] , \ab[16][17] ,
         \ab[16][16] , \ab[16][15] , \ab[16][14] , \ab[16][13] , \ab[16][12] ,
         \ab[16][11] , \ab[16][10] , \ab[16][9] , \ab[16][8] , \ab[16][7] ,
         \ab[16][6] , \ab[16][5] , \ab[16][4] , \ab[16][3] , \ab[16][2] ,
         \ab[16][1] , \ab[16][0] , \ab[15][31] , \ab[15][30] , \ab[15][29] ,
         \ab[15][28] , \ab[15][27] , \ab[15][26] , \ab[15][25] , \ab[15][24] ,
         \ab[15][23] , \ab[15][22] , \ab[15][21] , \ab[15][20] , \ab[15][19] ,
         \ab[15][18] , \ab[15][17] , \ab[15][16] , \ab[15][15] , \ab[15][14] ,
         \ab[15][13] , \ab[15][12] , \ab[15][11] , \ab[15][10] , \ab[15][9] ,
         \ab[15][8] , \ab[15][7] , \ab[15][6] , \ab[15][5] , \ab[15][4] ,
         \ab[15][3] , \ab[15][2] , \ab[15][1] , \ab[15][0] , \ab[14][31] ,
         \ab[14][30] , \ab[14][29] , \ab[14][28] , \ab[14][27] , \ab[14][26] ,
         \ab[14][25] , \ab[14][24] , \ab[14][23] , \ab[14][22] , \ab[14][21] ,
         \ab[14][20] , \ab[14][19] , \ab[14][18] , \ab[14][17] , \ab[14][16] ,
         \ab[14][15] , \ab[14][14] , \ab[14][13] , \ab[14][12] , \ab[14][11] ,
         \ab[14][10] , \ab[14][9] , \ab[14][8] , \ab[14][7] , \ab[14][6] ,
         \ab[14][5] , \ab[14][4] , \ab[14][3] , \ab[14][2] , \ab[14][1] ,
         \ab[14][0] , \ab[13][31] , \ab[13][30] , \ab[13][29] , \ab[13][28] ,
         \ab[13][27] , \ab[13][26] , \ab[13][25] , \ab[13][24] , \ab[13][23] ,
         \ab[13][22] , \ab[13][21] , \ab[13][20] , \ab[13][19] , \ab[13][18] ,
         \ab[13][17] , \ab[13][16] , \ab[13][15] , \ab[13][14] , \ab[13][13] ,
         \ab[13][12] , \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] ,
         \ab[13][7] , \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] ,
         \ab[13][2] , \ab[13][1] , \ab[13][0] , \ab[12][31] , \ab[12][30] ,
         \ab[12][29] , \ab[12][28] , \ab[12][27] , \ab[12][26] , \ab[12][25] ,
         \ab[12][24] , \ab[12][23] , \ab[12][22] , \ab[12][21] , \ab[12][20] ,
         \ab[12][19] , \ab[12][18] , \ab[12][17] , \ab[12][16] , \ab[12][15] ,
         \ab[12][14] , \ab[12][13] , \ab[12][12] , \ab[12][11] , \ab[12][10] ,
         \ab[12][9] , \ab[12][8] , \ab[12][7] , \ab[12][6] , \ab[12][5] ,
         \ab[12][4] , \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] ,
         \ab[11][31] , \ab[11][30] , \ab[11][29] , \ab[11][28] , \ab[11][27] ,
         \ab[11][26] , \ab[11][25] , \ab[11][24] , \ab[11][23] , \ab[11][22] ,
         \ab[11][21] , \ab[11][20] , \ab[11][19] , \ab[11][18] , \ab[11][17] ,
         \ab[11][16] , \ab[11][15] , \ab[11][14] , \ab[11][13] , \ab[11][12] ,
         \ab[11][11] , \ab[11][10] , \ab[11][9] , \ab[11][8] , \ab[11][7] ,
         \ab[11][6] , \ab[11][5] , \ab[11][4] , \ab[11][3] , \ab[11][2] ,
         \ab[11][1] , \ab[11][0] , \ab[10][31] , \ab[10][30] , \ab[10][29] ,
         \ab[10][28] , \ab[10][27] , \ab[10][26] , \ab[10][25] , \ab[10][24] ,
         \ab[10][23] , \ab[10][22] , \ab[10][21] , \ab[10][20] , \ab[10][19] ,
         \ab[10][18] , \ab[10][17] , \ab[10][16] , \ab[10][15] , \ab[10][14] ,
         \ab[10][13] , \ab[10][12] , \ab[10][11] , \ab[10][10] , \ab[10][9] ,
         \ab[10][8] , \ab[10][7] , \ab[10][6] , \ab[10][5] , \ab[10][4] ,
         \ab[10][3] , \ab[10][2] , \ab[10][1] , \ab[10][0] , \ab[9][31] ,
         \ab[9][30] , \ab[9][29] , \ab[9][28] , \ab[9][27] , \ab[9][26] ,
         \ab[9][25] , \ab[9][24] , \ab[9][23] , \ab[9][22] , \ab[9][21] ,
         \ab[9][20] , \ab[9][19] , \ab[9][18] , \ab[9][17] , \ab[9][16] ,
         \ab[9][15] , \ab[9][14] , \ab[9][13] , \ab[9][12] , \ab[9][11] ,
         \ab[9][10] , \ab[9][9] , \ab[9][8] , \ab[9][7] , \ab[9][6] ,
         \ab[9][5] , \ab[9][4] , \ab[9][3] , \ab[9][2] , \ab[9][1] ,
         \ab[9][0] , \ab[8][31] , \ab[8][30] , \ab[8][29] , \ab[8][28] ,
         \ab[8][27] , \ab[8][26] , \ab[8][25] , \ab[8][24] , \ab[8][23] ,
         \ab[8][22] , \ab[8][21] , \ab[8][20] , \ab[8][19] , \ab[8][18] ,
         \ab[8][17] , \ab[8][16] , \ab[8][15] , \ab[8][14] , \ab[8][13] ,
         \ab[8][12] , \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] ,
         \ab[8][7] , \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] ,
         \ab[8][2] , \ab[8][1] , \ab[8][0] , \ab[7][31] , \ab[7][30] ,
         \ab[7][29] , \ab[7][28] , \ab[7][27] , \ab[7][26] , \ab[7][25] ,
         \ab[7][24] , \ab[7][23] , \ab[7][22] , \ab[7][21] , \ab[7][20] ,
         \ab[7][19] , \ab[7][18] , \ab[7][17] , \ab[7][16] , \ab[7][15] ,
         \ab[7][14] , \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] ,
         \ab[7][9] , \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] ,
         \ab[7][4] , \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] ,
         \ab[6][31] , \ab[6][30] , \ab[6][29] , \ab[6][28] , \ab[6][27] ,
         \ab[6][26] , \ab[6][25] , \ab[6][24] , \ab[6][23] , \ab[6][22] ,
         \ab[6][21] , \ab[6][20] , \ab[6][19] , \ab[6][18] , \ab[6][17] ,
         \ab[6][16] , \ab[6][15] , \ab[6][14] , \ab[6][13] , \ab[6][12] ,
         \ab[6][11] , \ab[6][10] , \ab[6][9] , \ab[6][8] , \ab[6][7] ,
         \ab[6][6] , \ab[6][5] , \ab[6][4] , \ab[6][3] , \ab[6][2] ,
         \ab[6][1] , \ab[6][0] , \ab[5][31] , \ab[5][30] , \ab[5][29] ,
         \ab[5][28] , \ab[5][27] , \ab[5][26] , \ab[5][25] , \ab[5][24] ,
         \ab[5][23] , \ab[5][22] , \ab[5][21] , \ab[5][20] , \ab[5][19] ,
         \ab[5][18] , \ab[5][17] , \ab[5][16] , \ab[5][15] , \ab[5][14] ,
         \ab[5][13] , \ab[5][12] , \ab[5][11] , \ab[5][10] , \ab[5][9] ,
         \ab[5][8] , \ab[5][7] , \ab[5][6] , \ab[5][5] , \ab[5][4] ,
         \ab[5][3] , \ab[5][2] , \ab[5][1] , \ab[5][0] , \ab[4][31] ,
         \ab[4][30] , \ab[4][29] , \ab[4][28] , \ab[4][27] , \ab[4][26] ,
         \ab[4][25] , \ab[4][24] , \ab[4][23] , \ab[4][22] , \ab[4][21] ,
         \ab[4][20] , \ab[4][19] , \ab[4][18] , \ab[4][17] , \ab[4][16] ,
         \ab[4][15] , \ab[4][14] , \ab[4][13] , \ab[4][12] , \ab[4][11] ,
         \ab[4][10] , \ab[4][9] , \ab[4][8] , \ab[4][7] , \ab[4][6] ,
         \ab[4][5] , \ab[4][4] , \ab[4][3] , \ab[4][2] , \ab[4][1] ,
         \ab[4][0] , \ab[3][31] , \ab[3][30] , \ab[3][29] , \ab[3][28] ,
         \ab[3][27] , \ab[3][26] , \ab[3][25] , \ab[3][24] , \ab[3][23] ,
         \ab[3][22] , \ab[3][21] , \ab[3][20] , \ab[3][19] , \ab[3][18] ,
         \ab[3][17] , \ab[3][16] , \ab[3][15] , \ab[3][14] , \ab[3][13] ,
         \ab[3][12] , \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][8] ,
         \ab[3][7] , \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] ,
         \ab[3][2] , \ab[3][1] , \ab[3][0] , \ab[2][31] , \ab[2][30] ,
         \ab[2][29] , \ab[2][28] , \ab[2][27] , \ab[2][26] , \ab[2][25] ,
         \ab[2][24] , \ab[2][23] , \ab[2][22] , \ab[2][21] , \ab[2][20] ,
         \ab[2][19] , \ab[2][18] , \ab[2][17] , \ab[2][16] , \ab[2][15] ,
         \ab[2][14] , \ab[2][13] , \ab[2][12] , \ab[2][11] , \ab[2][10] ,
         \ab[2][9] , \ab[2][8] , \ab[2][7] , \ab[2][6] , \ab[2][5] ,
         \ab[2][4] , \ab[2][3] , \ab[2][2] , \ab[2][1] , \ab[2][0] ,
         \ab[1][31] , \ab[1][30] , \ab[1][29] , \ab[1][28] , \ab[1][27] ,
         \ab[1][26] , \ab[1][25] , \ab[1][24] , \ab[1][23] , \ab[1][22] ,
         \ab[1][21] , \ab[1][20] , \ab[1][19] , \ab[1][18] , \ab[1][17] ,
         \ab[1][16] , \ab[1][15] , \ab[1][14] , \ab[1][13] , \ab[1][12] ,
         \ab[1][11] , \ab[1][10] , \ab[1][9] , \ab[1][8] , \ab[1][7] ,
         \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] , \ab[1][2] ,
         \ab[1][1] , \ab[1][0] , \ab[0][31] , \ab[0][30] , \ab[0][29] ,
         \ab[0][28] , \ab[0][27] , \ab[0][26] , \ab[0][25] , \ab[0][24] ,
         \ab[0][23] , \ab[0][22] , \ab[0][21] , \ab[0][20] , \ab[0][19] ,
         \ab[0][18] , \ab[0][17] , \ab[0][16] , \ab[0][15] , \ab[0][14] ,
         \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] , \ab[0][9] ,
         \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] ,
         \ab[0][3] , \ab[0][2] , \ab[0][1] , \CARRYB[15][30] ,
         \CARRYB[15][29] , \CARRYB[15][28] , \CARRYB[15][27] ,
         \CARRYB[15][26] , \CARRYB[15][25] , \CARRYB[15][24] ,
         \CARRYB[15][23] , \CARRYB[15][22] , \CARRYB[15][21] ,
         \CARRYB[15][20] , \CARRYB[15][19] , \CARRYB[15][18] ,
         \CARRYB[15][17] , \CARRYB[15][16] , \CARRYB[15][15] ,
         \CARRYB[15][14] , \CARRYB[15][13] , \CARRYB[15][12] ,
         \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] ,
         \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] ,
         \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] ,
         \CARRYB[14][30] , \CARRYB[14][29] , \CARRYB[14][28] ,
         \CARRYB[14][27] , \CARRYB[14][26] , \CARRYB[14][25] ,
         \CARRYB[14][24] , \CARRYB[14][23] , \CARRYB[14][22] ,
         \CARRYB[14][21] , \CARRYB[14][20] , \CARRYB[14][19] ,
         \CARRYB[14][18] , \CARRYB[14][17] , \CARRYB[14][16] ,
         \CARRYB[14][15] , \CARRYB[14][14] , \CARRYB[14][13] ,
         \CARRYB[14][12] , \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] ,
         \CARRYB[14][8] , \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] ,
         \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] ,
         \CARRYB[14][0] , \CARRYB[13][30] , \CARRYB[13][29] , \CARRYB[13][28] ,
         \CARRYB[13][27] , \CARRYB[13][26] , \CARRYB[13][25] ,
         \CARRYB[13][24] , \CARRYB[13][23] , \CARRYB[13][22] ,
         \CARRYB[13][21] , \CARRYB[13][20] , \CARRYB[13][19] ,
         \CARRYB[13][18] , \CARRYB[13][17] , \CARRYB[13][16] ,
         \CARRYB[13][15] , \CARRYB[13][14] , \CARRYB[13][13] ,
         \CARRYB[13][12] , \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] ,
         \CARRYB[13][8] , \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] ,
         \CARRYB[13][4] , \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] ,
         \CARRYB[13][0] , \CARRYB[12][30] , \CARRYB[12][29] , \CARRYB[12][28] ,
         \CARRYB[12][27] , \CARRYB[12][26] , \CARRYB[12][25] ,
         \CARRYB[12][24] , \CARRYB[12][23] , \CARRYB[12][22] ,
         \CARRYB[12][21] , \CARRYB[12][20] , \CARRYB[12][19] ,
         \CARRYB[12][18] , \CARRYB[12][17] , \CARRYB[12][16] ,
         \CARRYB[12][15] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][30] , \CARRYB[11][29] , \CARRYB[11][28] ,
         \CARRYB[11][27] , \CARRYB[11][26] , \CARRYB[11][25] ,
         \CARRYB[11][24] , \CARRYB[11][23] , \CARRYB[11][22] ,
         \CARRYB[11][21] , \CARRYB[11][20] , \CARRYB[11][19] ,
         \CARRYB[11][18] , \CARRYB[11][17] , \CARRYB[11][16] ,
         \CARRYB[11][15] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][30] , \CARRYB[10][29] , \CARRYB[10][28] ,
         \CARRYB[10][27] , \CARRYB[10][26] , \CARRYB[10][25] ,
         \CARRYB[10][24] , \CARRYB[10][23] , \CARRYB[10][22] ,
         \CARRYB[10][21] , \CARRYB[10][20] , \CARRYB[10][19] ,
         \CARRYB[10][18] , \CARRYB[10][17] , \CARRYB[10][16] ,
         \CARRYB[10][15] , \CARRYB[10][14] , \CARRYB[10][13] ,
         \CARRYB[10][12] , \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] ,
         \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] ,
         \CARRYB[10][0] , \CARRYB[9][30] , \CARRYB[9][29] , \CARRYB[9][28] ,
         \CARRYB[9][27] , \CARRYB[9][26] , \CARRYB[9][25] , \CARRYB[9][24] ,
         \CARRYB[9][23] , \CARRYB[9][22] , \CARRYB[9][21] , \CARRYB[9][20] ,
         \CARRYB[9][19] , \CARRYB[9][18] , \CARRYB[9][17] , \CARRYB[9][16] ,
         \CARRYB[9][15] , \CARRYB[9][14] , \CARRYB[9][13] , \CARRYB[9][12] ,
         \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] , \CARRYB[9][8] ,
         \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][5] , \CARRYB[9][4] ,
         \CARRYB[9][3] , \CARRYB[9][2] , \CARRYB[9][1] , \CARRYB[9][0] ,
         \CARRYB[8][30] , \CARRYB[8][29] , \CARRYB[8][28] , \CARRYB[8][27] ,
         \CARRYB[8][26] , \CARRYB[8][25] , \CARRYB[8][24] , \CARRYB[8][23] ,
         \CARRYB[8][22] , \CARRYB[8][21] , \CARRYB[8][20] , \CARRYB[8][19] ,
         \CARRYB[8][18] , \CARRYB[8][17] , \CARRYB[8][16] , \CARRYB[8][15] ,
         \CARRYB[8][14] , \CARRYB[8][13] , \CARRYB[8][12] , \CARRYB[8][11] ,
         \CARRYB[8][10] , \CARRYB[8][9] , \CARRYB[8][8] , \CARRYB[8][7] ,
         \CARRYB[8][6] , \CARRYB[8][5] , \CARRYB[8][4] , \CARRYB[8][3] ,
         \CARRYB[8][2] , \CARRYB[8][1] , \CARRYB[8][0] , \CARRYB[7][30] ,
         \CARRYB[7][29] , \CARRYB[7][28] , \CARRYB[7][27] , \CARRYB[7][26] ,
         \CARRYB[7][25] , \CARRYB[7][24] , \CARRYB[7][23] , \CARRYB[7][22] ,
         \CARRYB[7][21] , \CARRYB[7][20] , \CARRYB[7][19] , \CARRYB[7][18] ,
         \CARRYB[7][17] , \CARRYB[7][16] , \CARRYB[7][15] , \CARRYB[7][14] ,
         \CARRYB[7][13] , \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] ,
         \CARRYB[7][9] , \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] ,
         \CARRYB[7][5] , \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] ,
         \CARRYB[7][1] , \CARRYB[7][0] , \CARRYB[6][30] , \CARRYB[6][29] ,
         \CARRYB[6][28] , \CARRYB[6][27] , \CARRYB[6][26] , \CARRYB[6][25] ,
         \CARRYB[6][24] , \CARRYB[6][23] , \CARRYB[6][22] , \CARRYB[6][21] ,
         \CARRYB[6][20] , \CARRYB[6][19] , \CARRYB[6][18] , \CARRYB[6][17] ,
         \CARRYB[6][16] , \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] ,
         \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] ,
         \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] ,
         \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][30] , \CARRYB[5][29] , \CARRYB[5][28] ,
         \CARRYB[5][27] , \CARRYB[5][26] , \CARRYB[5][25] , \CARRYB[5][24] ,
         \CARRYB[5][23] , \CARRYB[5][22] , \CARRYB[5][21] , \CARRYB[5][20] ,
         \CARRYB[5][19] , \CARRYB[5][18] , \CARRYB[5][17] , \CARRYB[5][16] ,
         \CARRYB[5][15] , \CARRYB[5][14] , \CARRYB[5][13] , \CARRYB[5][12] ,
         \CARRYB[5][11] , \CARRYB[5][10] , \CARRYB[5][9] , \CARRYB[5][8] ,
         \CARRYB[5][7] , \CARRYB[5][6] , \CARRYB[5][5] , \CARRYB[5][4] ,
         \CARRYB[5][3] , \CARRYB[5][2] , \CARRYB[5][1] , \CARRYB[5][0] ,
         \CARRYB[4][30] , \CARRYB[4][29] , \CARRYB[4][28] , \CARRYB[4][27] ,
         \CARRYB[4][26] , \CARRYB[4][25] , \CARRYB[4][24] , \CARRYB[4][23] ,
         \CARRYB[4][22] , \CARRYB[4][21] , \CARRYB[4][20] , \CARRYB[4][19] ,
         \CARRYB[4][18] , \CARRYB[4][17] , \CARRYB[4][16] , \CARRYB[4][15] ,
         \CARRYB[4][14] , \CARRYB[4][13] , \CARRYB[4][12] , \CARRYB[4][11] ,
         \CARRYB[4][10] , \CARRYB[4][9] , \CARRYB[4][8] , \CARRYB[4][7] ,
         \CARRYB[4][6] , \CARRYB[4][5] , \CARRYB[4][4] , \CARRYB[4][3] ,
         \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] , \CARRYB[3][30] ,
         \CARRYB[3][29] , \CARRYB[3][28] , \CARRYB[3][27] , \CARRYB[3][26] ,
         \CARRYB[3][25] , \CARRYB[3][24] , \CARRYB[3][23] , \CARRYB[3][22] ,
         \CARRYB[3][21] , \CARRYB[3][20] , \CARRYB[3][19] , \CARRYB[3][18] ,
         \CARRYB[3][17] , \CARRYB[3][16] , \CARRYB[3][15] , \CARRYB[3][14] ,
         \CARRYB[3][13] , \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] ,
         \CARRYB[3][9] , \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] ,
         \CARRYB[3][5] , \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] ,
         \CARRYB[3][1] , \CARRYB[3][0] , \CARRYB[2][30] , \CARRYB[2][29] ,
         \CARRYB[2][28] , \CARRYB[2][27] , \CARRYB[2][26] , \CARRYB[2][25] ,
         \CARRYB[2][24] , \CARRYB[2][23] , \CARRYB[2][22] , \CARRYB[2][21] ,
         \CARRYB[2][20] , \CARRYB[2][19] , \CARRYB[2][18] , \CARRYB[2][17] ,
         \CARRYB[2][16] , \CARRYB[2][15] , \CARRYB[2][14] , \CARRYB[2][13] ,
         \CARRYB[2][12] , \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] ,
         \CARRYB[2][8] , \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] ,
         \CARRYB[2][4] , \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] ,
         \CARRYB[2][0] , \CARRYB[1][30] , \CARRYB[1][29] , \CARRYB[1][28] ,
         \CARRYB[1][27] , \CARRYB[1][26] , \CARRYB[1][25] , \CARRYB[1][24] ,
         \CARRYB[1][23] , \CARRYB[1][22] , \CARRYB[1][21] , \CARRYB[1][20] ,
         \CARRYB[1][19] , \CARRYB[1][18] , \CARRYB[1][17] , \CARRYB[1][16] ,
         \CARRYB[1][15] , \CARRYB[1][14] , \CARRYB[1][13] , \CARRYB[1][12] ,
         \CARRYB[1][11] , \CARRYB[1][10] , \CARRYB[1][9] , \CARRYB[1][8] ,
         \CARRYB[1][7] , \CARRYB[1][6] , \CARRYB[1][5] , \CARRYB[1][4] ,
         \CARRYB[1][3] , \CARRYB[1][2] , \CARRYB[1][1] , \CARRYB[1][0] ,
         \SUMB[15][30] , \SUMB[15][29] , \SUMB[15][28] , \SUMB[15][27] ,
         \SUMB[15][26] , \SUMB[15][25] , \SUMB[15][24] , \SUMB[15][23] ,
         \SUMB[15][22] , \SUMB[15][21] , \SUMB[15][20] , \SUMB[15][19] ,
         \SUMB[15][18] , \SUMB[15][17] , \SUMB[15][16] , \SUMB[15][15] ,
         \SUMB[15][14] , \SUMB[15][13] , \SUMB[15][12] , \SUMB[15][11] ,
         \SUMB[15][10] , \SUMB[15][9] , \SUMB[15][8] , \SUMB[15][7] ,
         \SUMB[15][6] , \SUMB[15][5] , \SUMB[15][4] , \SUMB[15][3] ,
         \SUMB[15][2] , \SUMB[15][1] , \SUMB[14][30] , \SUMB[14][29] ,
         \SUMB[14][28] , \SUMB[14][27] , \SUMB[14][26] , \SUMB[14][25] ,
         \SUMB[14][24] , \SUMB[14][23] , \SUMB[14][22] , \SUMB[14][21] ,
         \SUMB[14][20] , \SUMB[14][19] , \SUMB[14][18] , \SUMB[14][17] ,
         \SUMB[14][16] , \SUMB[14][15] , \SUMB[14][14] , \SUMB[14][13] ,
         \SUMB[14][12] , \SUMB[14][11] , \SUMB[14][10] , \SUMB[14][9] ,
         \SUMB[14][8] , \SUMB[14][7] , \SUMB[14][6] , \SUMB[14][5] ,
         \SUMB[14][4] , \SUMB[14][3] , \SUMB[14][2] , \SUMB[14][1] ,
         \SUMB[13][30] , \SUMB[13][29] , \SUMB[13][28] , \SUMB[13][27] ,
         \SUMB[13][26] , \SUMB[13][25] , \SUMB[13][24] , \SUMB[13][23] ,
         \SUMB[13][22] , \SUMB[13][21] , \SUMB[13][20] , \SUMB[13][19] ,
         \SUMB[13][18] , \SUMB[13][17] , \SUMB[13][16] , \SUMB[13][15] ,
         \SUMB[13][14] , \SUMB[13][13] , \SUMB[13][12] , \SUMB[13][11] ,
         \SUMB[13][10] , \SUMB[13][9] , \SUMB[13][8] , \SUMB[13][7] ,
         \SUMB[13][6] , \SUMB[13][5] , \SUMB[13][4] , \SUMB[13][3] ,
         \SUMB[13][2] , \SUMB[13][1] , \SUMB[12][30] , \SUMB[12][29] ,
         \SUMB[12][28] , \SUMB[12][27] , \SUMB[12][26] , \SUMB[12][25] ,
         \SUMB[12][24] , \SUMB[12][23] , \SUMB[12][22] , \SUMB[12][21] ,
         \SUMB[12][20] , \SUMB[12][19] , \SUMB[12][18] , \SUMB[12][17] ,
         \SUMB[12][16] , \SUMB[12][15] , \SUMB[12][14] , \SUMB[12][13] ,
         \SUMB[12][12] , \SUMB[12][11] , \SUMB[12][10] , \SUMB[12][9] ,
         \SUMB[12][8] , \SUMB[12][7] , \SUMB[12][6] , \SUMB[12][5] ,
         \SUMB[12][4] , \SUMB[12][3] , \SUMB[12][2] , \SUMB[12][1] ,
         \SUMB[11][30] , \SUMB[11][29] , \SUMB[11][28] , \SUMB[11][27] ,
         \SUMB[11][26] , \SUMB[11][25] , \SUMB[11][24] , \SUMB[11][23] ,
         \SUMB[11][22] , \SUMB[11][21] , \SUMB[11][20] , \SUMB[11][19] ,
         \SUMB[11][18] , \SUMB[11][17] , \SUMB[11][16] , \SUMB[11][15] ,
         \SUMB[11][14] , \SUMB[11][13] , \SUMB[11][12] , \SUMB[11][11] ,
         \SUMB[11][10] , \SUMB[11][9] , \SUMB[11][8] , \SUMB[11][7] ,
         \SUMB[11][6] , \SUMB[11][5] , \SUMB[11][4] , \SUMB[11][3] ,
         \SUMB[11][2] , \SUMB[11][1] , \SUMB[10][30] , \SUMB[10][29] ,
         \SUMB[10][28] , \SUMB[10][27] , \SUMB[10][26] , \SUMB[10][25] ,
         \SUMB[10][24] , \SUMB[10][23] , \SUMB[10][22] , \SUMB[10][21] ,
         \SUMB[10][20] , \SUMB[10][19] , \SUMB[10][18] , \SUMB[10][17] ,
         \SUMB[10][16] , \SUMB[10][15] , \SUMB[10][14] , \SUMB[10][13] ,
         \SUMB[10][12] , \SUMB[10][11] , \SUMB[10][10] , \SUMB[10][9] ,
         \SUMB[10][8] , \SUMB[10][7] , \SUMB[10][6] , \SUMB[10][5] ,
         \SUMB[10][4] , \SUMB[10][3] , \SUMB[10][2] , \SUMB[10][1] ,
         \SUMB[9][30] , \SUMB[9][29] , \SUMB[9][28] , \SUMB[9][27] ,
         \SUMB[9][26] , \SUMB[9][25] , \SUMB[9][24] , \SUMB[9][23] ,
         \SUMB[9][22] , \SUMB[9][21] , \SUMB[9][20] , \SUMB[9][19] ,
         \SUMB[9][18] , \SUMB[9][17] , \SUMB[9][16] , \SUMB[9][15] ,
         \SUMB[9][14] , \SUMB[9][13] , \SUMB[9][12] , \SUMB[9][11] ,
         \SUMB[9][10] , \SUMB[9][9] , \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] ,
         \SUMB[9][5] , \SUMB[9][4] , \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] ,
         \SUMB[8][30] , \SUMB[8][29] , \SUMB[8][28] , \SUMB[8][27] ,
         \SUMB[8][26] , \SUMB[8][25] , \SUMB[8][24] , \SUMB[8][23] ,
         \SUMB[8][22] , \SUMB[8][21] , \SUMB[8][20] , \SUMB[8][19] ,
         \SUMB[8][18] , \SUMB[8][17] , \SUMB[8][16] , \SUMB[8][15] ,
         \SUMB[8][14] , \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] ,
         \SUMB[8][10] , \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] ,
         \SUMB[8][5] , \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] ,
         \SUMB[7][30] , \SUMB[7][29] , \SUMB[7][28] , \SUMB[7][27] ,
         \SUMB[7][26] , \SUMB[7][25] , \SUMB[7][24] , \SUMB[7][23] ,
         \SUMB[7][22] , \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] ,
         \SUMB[7][18] , \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] ,
         \SUMB[7][14] , \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] ,
         \SUMB[7][10] , \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] ,
         \SUMB[7][5] , \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] ,
         \SUMB[6][30] , \SUMB[6][29] , \SUMB[6][28] , \SUMB[6][27] ,
         \SUMB[6][26] , \SUMB[6][25] , \SUMB[6][24] , \SUMB[6][23] ,
         \SUMB[6][22] , \SUMB[6][21] , \SUMB[6][20] , \SUMB[6][19] ,
         \SUMB[6][18] , \SUMB[6][17] , \SUMB[6][16] , \SUMB[6][15] ,
         \SUMB[6][14] , \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] ,
         \SUMB[6][10] , \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] ,
         \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][30] , \SUMB[5][29] , \SUMB[5][28] , \SUMB[5][27] ,
         \SUMB[5][26] , \SUMB[5][25] , \SUMB[5][24] , \SUMB[5][23] ,
         \SUMB[5][22] , \SUMB[5][21] , \SUMB[5][20] , \SUMB[5][19] ,
         \SUMB[5][18] , \SUMB[5][17] , \SUMB[5][16] , \SUMB[5][15] ,
         \SUMB[5][14] , \SUMB[5][13] , \SUMB[5][12] , \SUMB[5][11] ,
         \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] , \SUMB[5][7] , \SUMB[5][6] ,
         \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] , \SUMB[5][2] , \SUMB[5][1] ,
         \SUMB[4][30] , \SUMB[4][29] , \SUMB[4][28] , \SUMB[4][27] ,
         \SUMB[4][26] , \SUMB[4][25] , \SUMB[4][24] , \SUMB[4][23] ,
         \SUMB[4][22] , \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] ,
         \SUMB[4][18] , \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] ,
         \SUMB[4][14] , \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] ,
         \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][30] , \SUMB[3][29] , \SUMB[3][28] , \SUMB[3][27] ,
         \SUMB[3][26] , \SUMB[3][25] , \SUMB[3][24] , \SUMB[3][23] ,
         \SUMB[3][22] , \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] ,
         \SUMB[3][18] , \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] ,
         \SUMB[3][14] , \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] ,
         \SUMB[3][10] , \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] ,
         \SUMB[3][5] , \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] ,
         \SUMB[2][30] , \SUMB[2][29] , \SUMB[2][28] , \SUMB[2][27] ,
         \SUMB[2][26] , \SUMB[2][25] , \SUMB[2][24] , \SUMB[2][23] ,
         \SUMB[2][22] , \SUMB[2][21] , \SUMB[2][20] , \SUMB[2][19] ,
         \SUMB[2][18] , \SUMB[2][17] , \SUMB[2][16] , \SUMB[2][15] ,
         \SUMB[2][14] , \SUMB[2][13] , \SUMB[2][12] , \SUMB[2][11] ,
         \SUMB[2][10] , \SUMB[2][9] , \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] ,
         \SUMB[2][5] , \SUMB[2][4] , \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] ,
         \SUMB[1][30] , \SUMB[1][29] , \SUMB[1][28] , \SUMB[1][27] ,
         \SUMB[1][26] , \SUMB[1][25] , \SUMB[1][24] , \SUMB[1][23] ,
         \SUMB[1][22] , \SUMB[1][21] , \SUMB[1][20] , \SUMB[1][19] ,
         \SUMB[1][18] , \SUMB[1][17] , \SUMB[1][16] , \SUMB[1][15] ,
         \SUMB[1][14] , \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] ,
         \SUMB[1][10] , \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] ,
         \SUMB[1][5] , \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] ,
         \CARRYB[31][31] , \CARRYB[31][30] , \CARRYB[31][29] ,
         \CARRYB[31][28] , \CARRYB[31][27] , \CARRYB[31][26] ,
         \CARRYB[31][25] , \CARRYB[31][24] , \CARRYB[31][23] ,
         \CARRYB[31][22] , \CARRYB[31][21] , \CARRYB[31][20] ,
         \CARRYB[31][19] , \CARRYB[31][18] , \CARRYB[31][17] ,
         \CARRYB[31][16] , \CARRYB[31][15] , \CARRYB[31][14] ,
         \CARRYB[31][13] , \CARRYB[31][12] , \CARRYB[31][11] ,
         \CARRYB[31][10] , \CARRYB[31][9] , \CARRYB[31][8] , \CARRYB[31][7] ,
         \CARRYB[31][6] , \CARRYB[31][5] , \CARRYB[31][4] , \CARRYB[31][3] ,
         \CARRYB[31][2] , \CARRYB[31][1] , \CARRYB[31][0] , \CARRYB[30][30] ,
         \CARRYB[30][29] , \CARRYB[30][28] , \CARRYB[30][27] ,
         \CARRYB[30][26] , \CARRYB[30][25] , \CARRYB[30][24] ,
         \CARRYB[30][23] , \CARRYB[30][22] , \CARRYB[30][21] ,
         \CARRYB[30][20] , \CARRYB[30][19] , \CARRYB[30][18] ,
         \CARRYB[30][17] , \CARRYB[30][16] , \CARRYB[30][15] ,
         \CARRYB[30][14] , \CARRYB[30][13] , \CARRYB[30][12] ,
         \CARRYB[30][11] , \CARRYB[30][10] , \CARRYB[30][9] , \CARRYB[30][8] ,
         \CARRYB[30][7] , \CARRYB[30][6] , \CARRYB[30][5] , \CARRYB[30][4] ,
         \CARRYB[30][3] , \CARRYB[30][2] , \CARRYB[30][1] , \CARRYB[30][0] ,
         \CARRYB[29][30] , \CARRYB[29][29] , \CARRYB[29][28] ,
         \CARRYB[29][27] , \CARRYB[29][26] , \CARRYB[29][25] ,
         \CARRYB[29][24] , \CARRYB[29][23] , \CARRYB[29][22] ,
         \CARRYB[29][21] , \CARRYB[29][20] , \CARRYB[29][19] ,
         \CARRYB[29][18] , \CARRYB[29][17] , \CARRYB[29][16] ,
         \CARRYB[29][15] , \CARRYB[29][14] , \CARRYB[29][13] ,
         \CARRYB[29][12] , \CARRYB[29][11] , \CARRYB[29][10] , \CARRYB[29][9] ,
         \CARRYB[29][8] , \CARRYB[29][7] , \CARRYB[29][6] , \CARRYB[29][5] ,
         \CARRYB[29][4] , \CARRYB[29][3] , \CARRYB[29][2] , \CARRYB[29][1] ,
         \CARRYB[29][0] , \CARRYB[28][30] , \CARRYB[28][29] , \CARRYB[28][28] ,
         \CARRYB[28][27] , \CARRYB[28][26] , \CARRYB[28][25] ,
         \CARRYB[28][24] , \CARRYB[28][23] , \CARRYB[28][22] ,
         \CARRYB[28][21] , \CARRYB[28][20] , \CARRYB[28][19] ,
         \CARRYB[28][18] , \CARRYB[28][17] , \CARRYB[28][16] ,
         \CARRYB[28][15] , \CARRYB[28][14] , \CARRYB[28][13] ,
         \CARRYB[28][12] , \CARRYB[28][11] , \CARRYB[28][10] , \CARRYB[28][9] ,
         \CARRYB[28][8] , \CARRYB[28][7] , \CARRYB[28][6] , \CARRYB[28][5] ,
         \CARRYB[28][4] , \CARRYB[28][3] , \CARRYB[28][2] , \CARRYB[28][1] ,
         \CARRYB[28][0] , \CARRYB[27][30] , \CARRYB[27][29] , \CARRYB[27][28] ,
         \CARRYB[27][27] , \CARRYB[27][26] , \CARRYB[27][25] ,
         \CARRYB[27][24] , \CARRYB[27][23] , \CARRYB[27][22] ,
         \CARRYB[27][21] , \CARRYB[27][20] , \CARRYB[27][19] ,
         \CARRYB[27][18] , \CARRYB[27][17] , \CARRYB[27][16] ,
         \CARRYB[27][15] , \CARRYB[27][14] , \CARRYB[27][13] ,
         \CARRYB[27][12] , \CARRYB[27][11] , \CARRYB[27][10] , \CARRYB[27][9] ,
         \CARRYB[27][8] , \CARRYB[27][7] , \CARRYB[27][6] , \CARRYB[27][5] ,
         \CARRYB[27][4] , \CARRYB[27][3] , \CARRYB[27][2] , \CARRYB[27][1] ,
         \CARRYB[27][0] , \CARRYB[26][30] , \CARRYB[26][29] , \CARRYB[26][28] ,
         \CARRYB[26][27] , \CARRYB[26][26] , \CARRYB[26][25] ,
         \CARRYB[26][24] , \CARRYB[26][23] , \CARRYB[26][22] ,
         \CARRYB[26][21] , \CARRYB[26][20] , \CARRYB[26][19] ,
         \CARRYB[26][18] , \CARRYB[26][17] , \CARRYB[26][16] ,
         \CARRYB[26][15] , \CARRYB[26][14] , \CARRYB[26][13] ,
         \CARRYB[26][12] , \CARRYB[26][11] , \CARRYB[26][10] , \CARRYB[26][9] ,
         \CARRYB[26][8] , \CARRYB[26][7] , \CARRYB[26][6] , \CARRYB[26][5] ,
         \CARRYB[26][4] , \CARRYB[26][3] , \CARRYB[26][2] , \CARRYB[26][1] ,
         \CARRYB[26][0] , \CARRYB[25][30] , \CARRYB[25][29] , \CARRYB[25][28] ,
         \CARRYB[25][27] , \CARRYB[25][26] , \CARRYB[25][25] ,
         \CARRYB[25][24] , \CARRYB[25][23] , \CARRYB[25][22] ,
         \CARRYB[25][21] , \CARRYB[25][20] , \CARRYB[25][19] ,
         \CARRYB[25][18] , \CARRYB[25][17] , \CARRYB[25][16] ,
         \CARRYB[25][15] , \CARRYB[25][14] , \CARRYB[25][13] ,
         \CARRYB[25][12] , \CARRYB[25][11] , \CARRYB[25][10] , \CARRYB[25][9] ,
         \CARRYB[25][8] , \CARRYB[25][7] , \CARRYB[25][6] , \CARRYB[25][5] ,
         \CARRYB[25][4] , \CARRYB[25][3] , \CARRYB[25][2] , \CARRYB[25][1] ,
         \CARRYB[25][0] , \CARRYB[24][30] , \CARRYB[24][29] , \CARRYB[24][28] ,
         \CARRYB[24][27] , \CARRYB[24][26] , \CARRYB[24][25] ,
         \CARRYB[24][24] , \CARRYB[24][23] , \CARRYB[24][22] ,
         \CARRYB[24][21] , \CARRYB[24][20] , \CARRYB[24][19] ,
         \CARRYB[24][18] , \CARRYB[24][17] , \CARRYB[24][16] ,
         \CARRYB[24][15] , \CARRYB[24][14] , \CARRYB[24][13] ,
         \CARRYB[24][12] , \CARRYB[24][11] , \CARRYB[24][10] , \CARRYB[24][9] ,
         \CARRYB[24][8] , \CARRYB[24][7] , \CARRYB[24][6] , \CARRYB[24][5] ,
         \CARRYB[24][4] , \CARRYB[24][3] , \CARRYB[24][2] , \CARRYB[24][1] ,
         \CARRYB[24][0] , \CARRYB[23][30] , \CARRYB[23][29] , \CARRYB[23][28] ,
         \CARRYB[23][27] , \CARRYB[23][26] , \CARRYB[23][25] ,
         \CARRYB[23][24] , \CARRYB[23][23] , \CARRYB[23][22] ,
         \CARRYB[23][21] , \CARRYB[23][20] , \CARRYB[23][19] ,
         \CARRYB[23][18] , \CARRYB[23][17] , \CARRYB[23][16] ,
         \CARRYB[23][15] , \CARRYB[23][14] , \CARRYB[23][13] ,
         \CARRYB[23][12] , \CARRYB[23][11] , \CARRYB[23][10] , \CARRYB[23][9] ,
         \CARRYB[23][8] , \CARRYB[23][7] , \CARRYB[23][6] , \CARRYB[23][5] ,
         \CARRYB[23][4] , \CARRYB[23][3] , \CARRYB[23][2] , \CARRYB[23][1] ,
         \CARRYB[23][0] , \CARRYB[22][30] , \CARRYB[22][29] , \CARRYB[22][28] ,
         \CARRYB[22][27] , \CARRYB[22][26] , \CARRYB[22][25] ,
         \CARRYB[22][24] , \CARRYB[22][23] , \CARRYB[22][22] ,
         \CARRYB[22][21] , \CARRYB[22][20] , \CARRYB[22][19] ,
         \CARRYB[22][18] , \CARRYB[22][17] , \CARRYB[22][16] ,
         \CARRYB[22][15] , \CARRYB[22][14] , \CARRYB[22][13] ,
         \CARRYB[22][12] , \CARRYB[22][11] , \CARRYB[22][10] , \CARRYB[22][9] ,
         \CARRYB[22][8] , \CARRYB[22][7] , \CARRYB[22][6] , \CARRYB[22][5] ,
         \CARRYB[22][4] , \CARRYB[22][3] , \CARRYB[22][2] , \CARRYB[22][1] ,
         \CARRYB[22][0] , \CARRYB[21][30] , \CARRYB[21][29] , \CARRYB[21][28] ,
         \CARRYB[21][27] , \CARRYB[21][26] , \CARRYB[21][25] ,
         \CARRYB[21][24] , \CARRYB[21][23] , \CARRYB[21][22] ,
         \CARRYB[21][21] , \CARRYB[21][20] , \CARRYB[21][19] ,
         \CARRYB[21][18] , \CARRYB[21][17] , \CARRYB[21][16] ,
         \CARRYB[21][15] , \CARRYB[21][14] , \CARRYB[21][13] ,
         \CARRYB[21][12] , \CARRYB[21][11] , \CARRYB[21][10] , \CARRYB[21][9] ,
         \CARRYB[21][8] , \CARRYB[21][7] , \CARRYB[21][6] , \CARRYB[21][5] ,
         \CARRYB[21][4] , \CARRYB[21][3] , \CARRYB[21][2] , \CARRYB[21][1] ,
         \CARRYB[21][0] , \CARRYB[20][30] , \CARRYB[20][29] , \CARRYB[20][28] ,
         \CARRYB[20][27] , \CARRYB[20][26] , \CARRYB[20][25] ,
         \CARRYB[20][24] , \CARRYB[20][23] , \CARRYB[20][22] ,
         \CARRYB[20][21] , \CARRYB[20][20] , \CARRYB[20][19] ,
         \CARRYB[20][18] , \CARRYB[20][17] , \CARRYB[20][16] ,
         \CARRYB[20][15] , \CARRYB[20][14] , \CARRYB[20][13] ,
         \CARRYB[20][12] , \CARRYB[20][11] , \CARRYB[20][10] , \CARRYB[20][9] ,
         \CARRYB[20][8] , \CARRYB[20][7] , \CARRYB[20][6] , \CARRYB[20][5] ,
         \CARRYB[20][4] , \CARRYB[20][3] , \CARRYB[20][2] , \CARRYB[20][1] ,
         \CARRYB[20][0] , \CARRYB[19][30] , \CARRYB[19][29] , \CARRYB[19][28] ,
         \CARRYB[19][27] , \CARRYB[19][26] , \CARRYB[19][25] ,
         \CARRYB[19][24] , \CARRYB[19][23] , \CARRYB[19][22] ,
         \CARRYB[19][21] , \CARRYB[19][20] , \CARRYB[19][19] ,
         \CARRYB[19][18] , \CARRYB[19][17] , \CARRYB[19][16] ,
         \CARRYB[19][15] , \CARRYB[19][14] , \CARRYB[19][13] ,
         \CARRYB[19][12] , \CARRYB[19][11] , \CARRYB[19][10] , \CARRYB[19][9] ,
         \CARRYB[19][8] , \CARRYB[19][7] , \CARRYB[19][6] , \CARRYB[19][5] ,
         \CARRYB[19][4] , \CARRYB[19][3] , \CARRYB[19][2] , \CARRYB[19][1] ,
         \CARRYB[19][0] , \CARRYB[18][30] , \CARRYB[18][29] , \CARRYB[18][28] ,
         \CARRYB[18][27] , \CARRYB[18][26] , \CARRYB[18][25] ,
         \CARRYB[18][24] , \CARRYB[18][23] , \CARRYB[18][22] ,
         \CARRYB[18][21] , \CARRYB[18][20] , \CARRYB[18][19] ,
         \CARRYB[18][18] , \CARRYB[18][17] , \CARRYB[18][16] ,
         \CARRYB[18][15] , \CARRYB[18][14] , \CARRYB[18][13] ,
         \CARRYB[18][12] , \CARRYB[18][11] , \CARRYB[18][10] , \CARRYB[18][9] ,
         \CARRYB[18][8] , \CARRYB[18][7] , \CARRYB[18][6] , \CARRYB[18][5] ,
         \CARRYB[18][4] , \CARRYB[18][3] , \CARRYB[18][2] , \CARRYB[18][1] ,
         \CARRYB[18][0] , \CARRYB[17][30] , \CARRYB[17][29] , \CARRYB[17][28] ,
         \CARRYB[17][27] , \CARRYB[17][26] , \CARRYB[17][25] ,
         \CARRYB[17][24] , \CARRYB[17][23] , \CARRYB[17][22] ,
         \CARRYB[17][21] , \CARRYB[17][20] , \CARRYB[17][19] ,
         \CARRYB[17][18] , \CARRYB[17][17] , \CARRYB[17][16] ,
         \CARRYB[17][15] , \CARRYB[17][14] , \CARRYB[17][13] ,
         \CARRYB[17][12] , \CARRYB[17][11] , \CARRYB[17][10] , \CARRYB[17][9] ,
         \CARRYB[17][8] , \CARRYB[17][7] , \CARRYB[17][6] , \CARRYB[17][5] ,
         \CARRYB[17][4] , \CARRYB[17][3] , \CARRYB[17][2] , \CARRYB[17][1] ,
         \CARRYB[17][0] , \CARRYB[16][30] , \CARRYB[16][29] , \CARRYB[16][28] ,
         \CARRYB[16][27] , \CARRYB[16][26] , \CARRYB[16][25] ,
         \CARRYB[16][24] , \CARRYB[16][23] , \CARRYB[16][22] ,
         \CARRYB[16][21] , \CARRYB[16][20] , \CARRYB[16][19] ,
         \CARRYB[16][18] , \CARRYB[16][17] , \CARRYB[16][16] ,
         \CARRYB[16][15] , \CARRYB[16][14] , \CARRYB[16][13] ,
         \CARRYB[16][12] , \CARRYB[16][11] , \CARRYB[16][10] , \CARRYB[16][9] ,
         \CARRYB[16][8] , \CARRYB[16][7] , \CARRYB[16][6] , \CARRYB[16][5] ,
         \CARRYB[16][4] , \CARRYB[16][3] , \CARRYB[16][2] , \CARRYB[16][1] ,
         \CARRYB[16][0] , \SUMB[31][31] , \SUMB[31][30] , \SUMB[31][29] ,
         \SUMB[31][28] , \SUMB[31][27] , \SUMB[31][26] , \SUMB[31][25] ,
         \SUMB[31][24] , \SUMB[31][23] , \SUMB[31][22] , \SUMB[31][21] ,
         \SUMB[31][20] , \SUMB[31][19] , \SUMB[31][18] , \SUMB[31][17] ,
         \SUMB[31][16] , \SUMB[31][15] , \SUMB[31][14] , \SUMB[31][13] ,
         \SUMB[31][12] , \SUMB[31][11] , \SUMB[31][10] , \SUMB[31][9] ,
         \SUMB[31][8] , \SUMB[31][7] , \SUMB[31][6] , \SUMB[31][5] ,
         \SUMB[31][4] , \SUMB[31][3] , \SUMB[31][2] , \SUMB[31][1] ,
         \SUMB[31][0] , \SUMB[30][30] , \SUMB[30][29] , \SUMB[30][28] ,
         \SUMB[30][27] , \SUMB[30][26] , \SUMB[30][25] , \SUMB[30][24] ,
         \SUMB[30][23] , \SUMB[30][22] , \SUMB[30][21] , \SUMB[30][20] ,
         \SUMB[30][19] , \SUMB[30][18] , \SUMB[30][17] , \SUMB[30][16] ,
         \SUMB[30][15] , \SUMB[30][14] , \SUMB[30][13] , \SUMB[30][12] ,
         \SUMB[30][11] , \SUMB[30][10] , \SUMB[30][9] , \SUMB[30][8] ,
         \SUMB[30][7] , \SUMB[30][6] , \SUMB[30][5] , \SUMB[30][4] ,
         \SUMB[30][3] , \SUMB[30][2] , \SUMB[30][1] , \SUMB[29][30] ,
         \SUMB[29][29] , \SUMB[29][28] , \SUMB[29][27] , \SUMB[29][26] ,
         \SUMB[29][25] , \SUMB[29][24] , \SUMB[29][23] , \SUMB[29][22] ,
         \SUMB[29][21] , \SUMB[29][20] , \SUMB[29][19] , \SUMB[29][18] ,
         \SUMB[29][17] , \SUMB[29][16] , \SUMB[29][15] , \SUMB[29][14] ,
         \SUMB[29][13] , \SUMB[29][12] , \SUMB[29][11] , \SUMB[29][10] ,
         \SUMB[29][9] , \SUMB[29][8] , \SUMB[29][7] , \SUMB[29][6] ,
         \SUMB[29][5] , \SUMB[29][4] , \SUMB[29][3] , \SUMB[29][2] ,
         \SUMB[29][1] , \SUMB[28][30] , \SUMB[28][29] , \SUMB[28][28] ,
         \SUMB[28][27] , \SUMB[28][26] , \SUMB[28][25] , \SUMB[28][24] ,
         \SUMB[28][23] , \SUMB[28][22] , \SUMB[28][21] , \SUMB[28][20] ,
         \SUMB[28][19] , \SUMB[28][18] , \SUMB[28][17] , \SUMB[28][16] ,
         \SUMB[28][15] , \SUMB[28][14] , \SUMB[28][13] , \SUMB[28][12] ,
         \SUMB[28][11] , \SUMB[28][10] , \SUMB[28][9] , \SUMB[28][8] ,
         \SUMB[28][7] , \SUMB[28][6] , \SUMB[28][5] , \SUMB[28][4] ,
         \SUMB[28][3] , \SUMB[28][2] , \SUMB[28][1] , \SUMB[27][30] ,
         \SUMB[27][29] , \SUMB[27][28] , \SUMB[27][27] , \SUMB[27][26] ,
         \SUMB[27][25] , \SUMB[27][24] , \SUMB[27][23] , \SUMB[27][22] ,
         \SUMB[27][21] , \SUMB[27][20] , \SUMB[27][19] , \SUMB[27][18] ,
         \SUMB[27][17] , \SUMB[27][16] , \SUMB[27][15] , \SUMB[27][14] ,
         \SUMB[27][13] , \SUMB[27][12] , \SUMB[27][11] , \SUMB[27][10] ,
         \SUMB[27][9] , \SUMB[27][8] , \SUMB[27][7] , \SUMB[27][6] ,
         \SUMB[27][5] , \SUMB[27][4] , \SUMB[27][3] , \SUMB[27][2] ,
         \SUMB[27][1] , \SUMB[26][30] , \SUMB[26][29] , \SUMB[26][28] ,
         \SUMB[26][27] , \SUMB[26][26] , \SUMB[26][25] , \SUMB[26][24] ,
         \SUMB[26][23] , \SUMB[26][22] , \SUMB[26][21] , \SUMB[26][20] ,
         \SUMB[26][19] , \SUMB[26][18] , \SUMB[26][17] , \SUMB[26][16] ,
         \SUMB[26][15] , \SUMB[26][14] , \SUMB[26][13] , \SUMB[26][12] ,
         \SUMB[26][11] , \SUMB[26][10] , \SUMB[26][9] , \SUMB[26][8] ,
         \SUMB[26][7] , \SUMB[26][6] , \SUMB[26][5] , \SUMB[26][4] ,
         \SUMB[26][3] , \SUMB[26][2] , \SUMB[26][1] , \SUMB[25][30] ,
         \SUMB[25][29] , \SUMB[25][28] , \SUMB[25][27] , \SUMB[25][26] ,
         \SUMB[25][25] , \SUMB[25][24] , \SUMB[25][23] , \SUMB[25][22] ,
         \SUMB[25][21] , \SUMB[25][20] , \SUMB[25][19] , \SUMB[25][18] ,
         \SUMB[25][17] , \SUMB[25][16] , \SUMB[25][15] , \SUMB[25][14] ,
         \SUMB[25][13] , \SUMB[25][12] , \SUMB[25][11] , \SUMB[25][10] ,
         \SUMB[25][9] , \SUMB[25][8] , \SUMB[25][7] , \SUMB[25][6] ,
         \SUMB[25][5] , \SUMB[25][4] , \SUMB[25][3] , \SUMB[25][2] ,
         \SUMB[25][1] , \SUMB[24][30] , \SUMB[24][29] , \SUMB[24][28] ,
         \SUMB[24][27] , \SUMB[24][26] , \SUMB[24][25] , \SUMB[24][24] ,
         \SUMB[24][23] , \SUMB[24][22] , \SUMB[24][21] , \SUMB[24][20] ,
         \SUMB[24][19] , \SUMB[24][18] , \SUMB[24][17] , \SUMB[24][16] ,
         \SUMB[24][15] , \SUMB[24][14] , \SUMB[24][13] , \SUMB[24][12] ,
         \SUMB[24][11] , \SUMB[24][10] , \SUMB[24][9] , \SUMB[24][8] ,
         \SUMB[24][7] , \SUMB[24][6] , \SUMB[24][5] , \SUMB[24][4] ,
         \SUMB[24][3] , \SUMB[24][2] , \SUMB[24][1] , \SUMB[23][30] ,
         \SUMB[23][29] , \SUMB[23][28] , \SUMB[23][27] , \SUMB[23][26] ,
         \SUMB[23][25] , \SUMB[23][24] , \SUMB[23][23] , \SUMB[23][22] ,
         \SUMB[23][21] , \SUMB[23][20] , \SUMB[23][19] , \SUMB[23][18] ,
         \SUMB[23][17] , \SUMB[23][16] , \SUMB[23][15] , \SUMB[23][14] ,
         \SUMB[23][13] , \SUMB[23][12] , \SUMB[23][11] , \SUMB[23][10] ,
         \SUMB[23][9] , \SUMB[23][8] , \SUMB[23][7] , \SUMB[23][6] ,
         \SUMB[23][5] , \SUMB[23][4] , \SUMB[23][3] , \SUMB[23][2] ,
         \SUMB[23][1] , \SUMB[22][30] , \SUMB[22][29] , \SUMB[22][28] ,
         \SUMB[22][27] , \SUMB[22][26] , \SUMB[22][25] , \SUMB[22][24] ,
         \SUMB[22][23] , \SUMB[22][22] , \SUMB[22][21] , \SUMB[22][20] ,
         \SUMB[22][19] , \SUMB[22][18] , \SUMB[22][17] , \SUMB[22][16] ,
         \SUMB[22][15] , \SUMB[22][14] , \SUMB[22][13] , \SUMB[22][12] ,
         \SUMB[22][11] , \SUMB[22][10] , \SUMB[22][9] , \SUMB[22][8] ,
         \SUMB[22][7] , \SUMB[22][6] , \SUMB[22][5] , \SUMB[22][4] ,
         \SUMB[22][3] , \SUMB[22][2] , \SUMB[22][1] , \SUMB[21][30] ,
         \SUMB[21][29] , \SUMB[21][28] , \SUMB[21][27] , \SUMB[21][26] ,
         \SUMB[21][25] , \SUMB[21][24] , \SUMB[21][23] , \SUMB[21][22] ,
         \SUMB[21][21] , \SUMB[21][20] , \SUMB[21][19] , \SUMB[21][18] ,
         \SUMB[21][17] , \SUMB[21][16] , \SUMB[21][15] , \SUMB[21][14] ,
         \SUMB[21][13] , \SUMB[21][12] , \SUMB[21][11] , \SUMB[21][10] ,
         \SUMB[21][9] , \SUMB[21][8] , \SUMB[21][7] , \SUMB[21][6] ,
         \SUMB[21][5] , \SUMB[21][4] , \SUMB[21][3] , \SUMB[21][2] ,
         \SUMB[21][1] , \SUMB[20][30] , \SUMB[20][29] , \SUMB[20][28] ,
         \SUMB[20][27] , \SUMB[20][26] , \SUMB[20][25] , \SUMB[20][24] ,
         \SUMB[20][23] , \SUMB[20][22] , \SUMB[20][21] , \SUMB[20][20] ,
         \SUMB[20][19] , \SUMB[20][18] , \SUMB[20][17] , \SUMB[20][16] ,
         \SUMB[20][15] , \SUMB[20][14] , \SUMB[20][13] , \SUMB[20][12] ,
         \SUMB[20][11] , \SUMB[20][10] , \SUMB[20][9] , \SUMB[20][8] ,
         \SUMB[20][7] , \SUMB[20][6] , \SUMB[20][5] , \SUMB[20][4] ,
         \SUMB[20][3] , \SUMB[20][2] , \SUMB[20][1] , \SUMB[19][30] ,
         \SUMB[19][29] , \SUMB[19][28] , \SUMB[19][27] , \SUMB[19][26] ,
         \SUMB[19][25] , \SUMB[19][24] , \SUMB[19][23] , \SUMB[19][22] ,
         \SUMB[19][21] , \SUMB[19][20] , \SUMB[19][19] , \SUMB[19][18] ,
         \SUMB[19][17] , \SUMB[19][16] , \SUMB[19][15] , \SUMB[19][14] ,
         \SUMB[19][13] , \SUMB[19][12] , \SUMB[19][11] , \SUMB[19][10] ,
         \SUMB[19][9] , \SUMB[19][8] , \SUMB[19][7] , \SUMB[19][6] ,
         \SUMB[19][5] , \SUMB[19][4] , \SUMB[19][3] , \SUMB[19][2] ,
         \SUMB[19][1] , \SUMB[18][30] , \SUMB[18][29] , \SUMB[18][28] ,
         \SUMB[18][27] , \SUMB[18][26] , \SUMB[18][25] , \SUMB[18][24] ,
         \SUMB[18][23] , \SUMB[18][22] , \SUMB[18][21] , \SUMB[18][20] ,
         \SUMB[18][19] , \SUMB[18][18] , \SUMB[18][17] , \SUMB[18][16] ,
         \SUMB[18][15] , \SUMB[18][14] , \SUMB[18][13] , \SUMB[18][12] ,
         \SUMB[18][11] , \SUMB[18][10] , \SUMB[18][9] , \SUMB[18][8] ,
         \SUMB[18][7] , \SUMB[18][6] , \SUMB[18][5] , \SUMB[18][4] ,
         \SUMB[18][3] , \SUMB[18][2] , \SUMB[18][1] , \SUMB[17][30] ,
         \SUMB[17][29] , \SUMB[17][28] , \SUMB[17][27] , \SUMB[17][26] ,
         \SUMB[17][25] , \SUMB[17][24] , \SUMB[17][23] , \SUMB[17][22] ,
         \SUMB[17][21] , \SUMB[17][20] , \SUMB[17][19] , \SUMB[17][18] ,
         \SUMB[17][17] , \SUMB[17][16] , \SUMB[17][15] , \SUMB[17][14] ,
         \SUMB[17][13] , \SUMB[17][12] , \SUMB[17][11] , \SUMB[17][10] ,
         \SUMB[17][9] , \SUMB[17][8] , \SUMB[17][7] , \SUMB[17][6] ,
         \SUMB[17][5] , \SUMB[17][4] , \SUMB[17][3] , \SUMB[17][2] ,
         \SUMB[17][1] , \SUMB[16][30] , \SUMB[16][29] , \SUMB[16][28] ,
         \SUMB[16][27] , \SUMB[16][26] , \SUMB[16][25] , \SUMB[16][24] ,
         \SUMB[16][23] , \SUMB[16][22] , \SUMB[16][21] , \SUMB[16][20] ,
         \SUMB[16][19] , \SUMB[16][18] , \SUMB[16][17] , \SUMB[16][16] ,
         \SUMB[16][15] , \SUMB[16][14] , \SUMB[16][13] , \SUMB[16][12] ,
         \SUMB[16][11] , \SUMB[16][10] , \SUMB[16][9] , \SUMB[16][8] ,
         \SUMB[16][7] , \SUMB[16][6] , \SUMB[16][5] , \SUMB[16][4] ,
         \SUMB[16][3] , \SUMB[16][2] , \SUMB[16][1] , QA, QB, ZA, ZB, \A1[61] ,
         \A1[60] , \A1[59] , \A1[58] , \A1[57] , \A1[56] , \A1[55] , \A1[54] ,
         \A1[53] , \A1[52] , \A1[51] , \A1[50] , \A1[49] , \A1[48] , \A1[47] ,
         \A1[46] , \A1[45] , \A1[44] , \A1[43] , \A1[42] , \A1[41] , \A1[40] ,
         \A1[39] , \A1[38] , \A1[37] , \A1[36] , \A1[35] , \A1[34] , \A1[33] ,
         \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] , \A1[27] , \A1[26] ,
         \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] ,
         \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] ,
         \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] ,
         \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] , \A2[61] , \A2[60] ,
         \A2[59] , \A2[58] , \A2[57] , \A2[56] , \A2[55] , \A2[54] , \A2[53] ,
         \A2[52] , \A2[51] , \A2[50] , \A2[49] , \A2[48] , \A2[47] , \A2[46] ,
         \A2[45] , \A2[44] , \A2[43] , \A2[42] , \A2[41] , \A2[40] , \A2[39] ,
         \A2[38] , \A2[37] , \A2[36] , \A2[35] , \A2[34] , \A2[33] , \A2[32] ,
         \A2[31] , \A2[30] , n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12,
         n13, n14, n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n66, n67, n68, n69, n70,
         n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84,
         n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98,
         n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109, n110,
         n111, n112, n113, n114, n115, n116, n117, n118, n119, n120, n121,
         n122, n123, n124, n125, n126, n127, n128, n129, n130, n131, n132,
         n133, n134, n135, n136, n137, n138, n139, n140, n141, n142, n143,
         n144, n145, n146, n147, n148, n149, n150, n151, n152, n153, n154,
         n155, n156, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n166, n167, n168, n169, n170, n171, n172, n173, n174, n175, n176,
         n177, n178, n179, n180, n181, n182, n183, n184, n185, n186, n187,
         n188, n189, n190, n191, n192, n193, n194, n195, n196, n197, n198,
         n199, n200, n201, n202, n203, n204, n205, n206, n207, n208, n209,
         n210;
  assign ZA = A[31];
  assign ZB = B[31];

  FA_X1 S14_31_0 ( .A(ZA), .B(ZB), .CI(\SUMB[31][0] ), .CO(\A2[30] ), .S(
        \A1[29] ) );
  FA_X1 S4_0 ( .A(\ab[31][0] ), .B(\CARRYB[30][0] ), .CI(\SUMB[30][1] ), .CO(
        \CARRYB[31][0] ), .S(\SUMB[31][0] ) );
  FA_X1 S4_2 ( .A(\ab[31][2] ), .B(\CARRYB[30][2] ), .CI(\SUMB[30][3] ), .CO(
        \CARRYB[31][2] ), .S(\SUMB[31][2] ) );
  FA_X1 S4_3 ( .A(\CARRYB[30][3] ), .B(\ab[31][3] ), .CI(\SUMB[30][4] ), .CO(
        \CARRYB[31][3] ), .S(\SUMB[31][3] ) );
  FA_X1 S4_4 ( .A(\CARRYB[30][4] ), .B(\ab[31][4] ), .CI(\SUMB[30][5] ), .CO(
        \CARRYB[31][4] ), .S(\SUMB[31][4] ) );
  FA_X1 S4_5 ( .A(\ab[31][5] ), .B(\CARRYB[30][5] ), .CI(\SUMB[30][6] ), .CO(
        \CARRYB[31][5] ), .S(\SUMB[31][5] ) );
  FA_X1 S4_6 ( .A(\ab[31][6] ), .B(\CARRYB[30][6] ), .CI(\SUMB[30][7] ), .CO(
        \CARRYB[31][6] ), .S(\SUMB[31][6] ) );
  FA_X1 S4_7 ( .A(\ab[31][7] ), .B(\CARRYB[30][7] ), .CI(\SUMB[30][8] ), .CO(
        \CARRYB[31][7] ), .S(\SUMB[31][7] ) );
  FA_X1 S4_8 ( .A(\ab[31][8] ), .B(\CARRYB[30][8] ), .CI(\SUMB[30][9] ), .CO(
        \CARRYB[31][8] ), .S(\SUMB[31][8] ) );
  FA_X1 S4_9 ( .A(\ab[31][9] ), .B(\CARRYB[30][9] ), .CI(\SUMB[30][10] ), .CO(
        \CARRYB[31][9] ), .S(\SUMB[31][9] ) );
  FA_X1 S4_10 ( .A(\ab[31][10] ), .B(\CARRYB[30][10] ), .CI(\SUMB[30][11] ), 
        .CO(\CARRYB[31][10] ), .S(\SUMB[31][10] ) );
  FA_X1 S4_11 ( .A(\ab[31][11] ), .B(\CARRYB[30][11] ), .CI(\SUMB[30][12] ), 
        .CO(\CARRYB[31][11] ), .S(\SUMB[31][11] ) );
  FA_X1 S4_12 ( .A(\ab[31][12] ), .B(\CARRYB[30][12] ), .CI(\SUMB[30][13] ), 
        .CO(\CARRYB[31][12] ), .S(\SUMB[31][12] ) );
  FA_X1 S4_13 ( .A(\ab[31][13] ), .B(\CARRYB[30][13] ), .CI(\SUMB[30][14] ), 
        .CO(\CARRYB[31][13] ), .S(\SUMB[31][13] ) );
  FA_X1 S4_14 ( .A(\ab[31][14] ), .B(\CARRYB[30][14] ), .CI(\SUMB[30][15] ), 
        .CO(\CARRYB[31][14] ), .S(\SUMB[31][14] ) );
  FA_X1 S4_15 ( .A(\ab[31][15] ), .B(\CARRYB[30][15] ), .CI(\SUMB[30][16] ), 
        .CO(\CARRYB[31][15] ), .S(\SUMB[31][15] ) );
  FA_X1 S4_16 ( .A(\ab[31][16] ), .B(\CARRYB[30][16] ), .CI(\SUMB[30][17] ), 
        .CO(\CARRYB[31][16] ), .S(\SUMB[31][16] ) );
  FA_X1 S4_17 ( .A(\ab[31][17] ), .B(\CARRYB[30][17] ), .CI(\SUMB[30][18] ), 
        .CO(\CARRYB[31][17] ), .S(\SUMB[31][17] ) );
  FA_X1 S4_18 ( .A(\ab[31][18] ), .B(\CARRYB[30][18] ), .CI(\SUMB[30][19] ), 
        .CO(\CARRYB[31][18] ), .S(\SUMB[31][18] ) );
  FA_X1 S4_19 ( .A(\ab[31][19] ), .B(\CARRYB[30][19] ), .CI(\SUMB[30][20] ), 
        .CO(\CARRYB[31][19] ), .S(\SUMB[31][19] ) );
  FA_X1 S4_20 ( .A(\ab[31][20] ), .B(\CARRYB[30][20] ), .CI(\SUMB[30][21] ), 
        .CO(\CARRYB[31][20] ), .S(\SUMB[31][20] ) );
  FA_X1 S4_21 ( .A(\ab[31][21] ), .B(\CARRYB[30][21] ), .CI(\SUMB[30][22] ), 
        .CO(\CARRYB[31][21] ), .S(\SUMB[31][21] ) );
  FA_X1 S4_22 ( .A(\ab[31][22] ), .B(\CARRYB[30][22] ), .CI(\SUMB[30][23] ), 
        .CO(\CARRYB[31][22] ), .S(\SUMB[31][22] ) );
  FA_X1 S4_23 ( .A(\ab[31][23] ), .B(\CARRYB[30][23] ), .CI(\SUMB[30][24] ), 
        .CO(\CARRYB[31][23] ), .S(\SUMB[31][23] ) );
  FA_X1 S4_24 ( .A(\ab[31][24] ), .B(\CARRYB[30][24] ), .CI(\SUMB[30][25] ), 
        .CO(\CARRYB[31][24] ), .S(\SUMB[31][24] ) );
  FA_X1 S4_25 ( .A(\ab[31][25] ), .B(\CARRYB[30][25] ), .CI(\SUMB[30][26] ), 
        .CO(\CARRYB[31][25] ), .S(\SUMB[31][25] ) );
  FA_X1 S4_26 ( .A(\ab[31][26] ), .B(\CARRYB[30][26] ), .CI(\SUMB[30][27] ), 
        .CO(\CARRYB[31][26] ), .S(\SUMB[31][26] ) );
  FA_X1 S4_27 ( .A(\ab[31][27] ), .B(\CARRYB[30][27] ), .CI(\SUMB[30][28] ), 
        .CO(\CARRYB[31][27] ), .S(\SUMB[31][27] ) );
  FA_X1 S4_28 ( .A(\ab[31][28] ), .B(\CARRYB[30][28] ), .CI(\SUMB[30][29] ), 
        .CO(\CARRYB[31][28] ), .S(\SUMB[31][28] ) );
  FA_X1 S4_29 ( .A(\ab[31][29] ), .B(\CARRYB[30][29] ), .CI(\SUMB[30][30] ), 
        .CO(\CARRYB[31][29] ), .S(\SUMB[31][29] ) );
  FA_X1 S5_30 ( .A(\ab[31][30] ), .B(\CARRYB[30][30] ), .CI(\ab[30][31] ), 
        .CO(\CARRYB[31][30] ), .S(\SUMB[31][30] ) );
  FA_X1 S14_31 ( .A(n210), .B(n208), .CI(\ab[31][31] ), .CO(\CARRYB[31][31] ), 
        .S(\SUMB[31][31] ) );
  FA_X1 S1_30_0 ( .A(\ab[30][0] ), .B(\CARRYB[29][0] ), .CI(\SUMB[29][1] ), 
        .CO(\CARRYB[30][0] ), .S(\A1[28] ) );
  FA_X1 S2_30_1 ( .A(\CARRYB[29][1] ), .B(\ab[30][1] ), .CI(\SUMB[29][2] ), 
        .CO(\CARRYB[30][1] ), .S(\SUMB[30][1] ) );
  FA_X1 S2_30_2 ( .A(\ab[30][2] ), .B(\CARRYB[29][2] ), .CI(\SUMB[29][3] ), 
        .CO(\CARRYB[30][2] ), .S(\SUMB[30][2] ) );
  FA_X1 S2_30_3 ( .A(\ab[30][3] ), .B(\CARRYB[29][3] ), .CI(\SUMB[29][4] ), 
        .CO(\CARRYB[30][3] ), .S(\SUMB[30][3] ) );
  FA_X1 S2_30_4 ( .A(\CARRYB[29][4] ), .B(\ab[30][4] ), .CI(\SUMB[29][5] ), 
        .CO(\CARRYB[30][4] ), .S(\SUMB[30][4] ) );
  FA_X1 S2_30_5 ( .A(\CARRYB[29][5] ), .B(\ab[30][5] ), .CI(\SUMB[29][6] ), 
        .CO(\CARRYB[30][5] ), .S(\SUMB[30][5] ) );
  FA_X1 S2_30_6 ( .A(\ab[30][6] ), .B(\CARRYB[29][6] ), .CI(\SUMB[29][7] ), 
        .CO(\CARRYB[30][6] ), .S(\SUMB[30][6] ) );
  FA_X1 S2_30_7 ( .A(\ab[30][7] ), .B(\CARRYB[29][7] ), .CI(\SUMB[29][8] ), 
        .CO(\CARRYB[30][7] ), .S(\SUMB[30][7] ) );
  FA_X1 S2_30_8 ( .A(\ab[30][8] ), .B(\CARRYB[29][8] ), .CI(\SUMB[29][9] ), 
        .CO(\CARRYB[30][8] ), .S(\SUMB[30][8] ) );
  FA_X1 S2_30_9 ( .A(\ab[30][9] ), .B(\CARRYB[29][9] ), .CI(\SUMB[29][10] ), 
        .CO(\CARRYB[30][9] ), .S(\SUMB[30][9] ) );
  FA_X1 S2_30_10 ( .A(\ab[30][10] ), .B(\CARRYB[29][10] ), .CI(\SUMB[29][11] ), 
        .CO(\CARRYB[30][10] ), .S(\SUMB[30][10] ) );
  FA_X1 S2_30_11 ( .A(\ab[30][11] ), .B(\CARRYB[29][11] ), .CI(\SUMB[29][12] ), 
        .CO(\CARRYB[30][11] ), .S(\SUMB[30][11] ) );
  FA_X1 S2_30_12 ( .A(\ab[30][12] ), .B(\CARRYB[29][12] ), .CI(\SUMB[29][13] ), 
        .CO(\CARRYB[30][12] ), .S(\SUMB[30][12] ) );
  FA_X1 S2_30_13 ( .A(\ab[30][13] ), .B(\CARRYB[29][13] ), .CI(\SUMB[29][14] ), 
        .CO(\CARRYB[30][13] ), .S(\SUMB[30][13] ) );
  FA_X1 S2_30_14 ( .A(\ab[30][14] ), .B(\CARRYB[29][14] ), .CI(\SUMB[29][15] ), 
        .CO(\CARRYB[30][14] ), .S(\SUMB[30][14] ) );
  FA_X1 S2_30_15 ( .A(\ab[30][15] ), .B(\CARRYB[29][15] ), .CI(\SUMB[29][16] ), 
        .CO(\CARRYB[30][15] ), .S(\SUMB[30][15] ) );
  FA_X1 S2_30_16 ( .A(\ab[30][16] ), .B(\CARRYB[29][16] ), .CI(\SUMB[29][17] ), 
        .CO(\CARRYB[30][16] ), .S(\SUMB[30][16] ) );
  FA_X1 S2_30_17 ( .A(\ab[30][17] ), .B(\CARRYB[29][17] ), .CI(\SUMB[29][18] ), 
        .CO(\CARRYB[30][17] ), .S(\SUMB[30][17] ) );
  FA_X1 S2_30_18 ( .A(\ab[30][18] ), .B(\CARRYB[29][18] ), .CI(\SUMB[29][19] ), 
        .CO(\CARRYB[30][18] ), .S(\SUMB[30][18] ) );
  FA_X1 S2_30_19 ( .A(\ab[30][19] ), .B(\CARRYB[29][19] ), .CI(\SUMB[29][20] ), 
        .CO(\CARRYB[30][19] ), .S(\SUMB[30][19] ) );
  FA_X1 S2_30_20 ( .A(\ab[30][20] ), .B(\CARRYB[29][20] ), .CI(\SUMB[29][21] ), 
        .CO(\CARRYB[30][20] ), .S(\SUMB[30][20] ) );
  FA_X1 S2_30_21 ( .A(\ab[30][21] ), .B(\CARRYB[29][21] ), .CI(\SUMB[29][22] ), 
        .CO(\CARRYB[30][21] ), .S(\SUMB[30][21] ) );
  FA_X1 S2_30_22 ( .A(\ab[30][22] ), .B(\CARRYB[29][22] ), .CI(\SUMB[29][23] ), 
        .CO(\CARRYB[30][22] ), .S(\SUMB[30][22] ) );
  FA_X1 S2_30_23 ( .A(\ab[30][23] ), .B(\CARRYB[29][23] ), .CI(\SUMB[29][24] ), 
        .CO(\CARRYB[30][23] ), .S(\SUMB[30][23] ) );
  FA_X1 S2_30_24 ( .A(\ab[30][24] ), .B(\CARRYB[29][24] ), .CI(\SUMB[29][25] ), 
        .CO(\CARRYB[30][24] ), .S(\SUMB[30][24] ) );
  FA_X1 S2_30_25 ( .A(\ab[30][25] ), .B(\CARRYB[29][25] ), .CI(\SUMB[29][26] ), 
        .CO(\CARRYB[30][25] ), .S(\SUMB[30][25] ) );
  FA_X1 S2_30_26 ( .A(\ab[30][26] ), .B(\CARRYB[29][26] ), .CI(\SUMB[29][27] ), 
        .CO(\CARRYB[30][26] ), .S(\SUMB[30][26] ) );
  FA_X1 S2_30_27 ( .A(\ab[30][27] ), .B(\CARRYB[29][27] ), .CI(\SUMB[29][28] ), 
        .CO(\CARRYB[30][27] ), .S(\SUMB[30][27] ) );
  FA_X1 S2_30_28 ( .A(\ab[30][28] ), .B(\CARRYB[29][28] ), .CI(\SUMB[29][29] ), 
        .CO(\CARRYB[30][28] ), .S(\SUMB[30][28] ) );
  FA_X1 S2_30_29 ( .A(\ab[30][29] ), .B(\CARRYB[29][29] ), .CI(\SUMB[29][30] ), 
        .CO(\CARRYB[30][29] ), .S(\SUMB[30][29] ) );
  FA_X1 S3_30_30 ( .A(\ab[30][30] ), .B(\CARRYB[29][30] ), .CI(\ab[29][31] ), 
        .CO(\CARRYB[30][30] ), .S(\SUMB[30][30] ) );
  FA_X1 S1_29_0 ( .A(\ab[29][0] ), .B(\CARRYB[28][0] ), .CI(\SUMB[28][1] ), 
        .CO(\CARRYB[29][0] ), .S(\A1[27] ) );
  FA_X1 S2_29_1 ( .A(\ab[29][1] ), .B(\CARRYB[28][1] ), .CI(\SUMB[28][2] ), 
        .CO(\CARRYB[29][1] ), .S(\SUMB[29][1] ) );
  FA_X1 S2_29_2 ( .A(\ab[29][2] ), .B(\CARRYB[28][2] ), .CI(\SUMB[28][3] ), 
        .CO(\CARRYB[29][2] ), .S(\SUMB[29][2] ) );
  FA_X1 S2_29_3 ( .A(\ab[29][3] ), .B(\CARRYB[28][3] ), .CI(\SUMB[28][4] ), 
        .CO(\CARRYB[29][3] ), .S(\SUMB[29][3] ) );
  FA_X1 S2_29_4 ( .A(\ab[29][4] ), .B(\CARRYB[28][4] ), .CI(\SUMB[28][5] ), 
        .CO(\CARRYB[29][4] ), .S(\SUMB[29][4] ) );
  FA_X1 S2_29_5 ( .A(\CARRYB[28][5] ), .B(\ab[29][5] ), .CI(\SUMB[28][6] ), 
        .CO(\CARRYB[29][5] ), .S(\SUMB[29][5] ) );
  FA_X1 S2_29_6 ( .A(\ab[29][6] ), .B(\CARRYB[28][6] ), .CI(\SUMB[28][7] ), 
        .CO(\CARRYB[29][6] ), .S(\SUMB[29][6] ) );
  FA_X1 S2_29_7 ( .A(\ab[29][7] ), .B(\CARRYB[28][7] ), .CI(\SUMB[28][8] ), 
        .CO(\CARRYB[29][7] ), .S(\SUMB[29][7] ) );
  FA_X1 S2_29_8 ( .A(\ab[29][8] ), .B(\CARRYB[28][8] ), .CI(\SUMB[28][9] ), 
        .CO(\CARRYB[29][8] ), .S(\SUMB[29][8] ) );
  FA_X1 S2_29_9 ( .A(\ab[29][9] ), .B(\CARRYB[28][9] ), .CI(\SUMB[28][10] ), 
        .CO(\CARRYB[29][9] ), .S(\SUMB[29][9] ) );
  FA_X1 S2_29_10 ( .A(\ab[29][10] ), .B(\CARRYB[28][10] ), .CI(\SUMB[28][11] ), 
        .CO(\CARRYB[29][10] ), .S(\SUMB[29][10] ) );
  FA_X1 S2_29_11 ( .A(\ab[29][11] ), .B(\CARRYB[28][11] ), .CI(\SUMB[28][12] ), 
        .CO(\CARRYB[29][11] ), .S(\SUMB[29][11] ) );
  FA_X1 S2_29_12 ( .A(\ab[29][12] ), .B(\CARRYB[28][12] ), .CI(\SUMB[28][13] ), 
        .CO(\CARRYB[29][12] ), .S(\SUMB[29][12] ) );
  FA_X1 S2_29_13 ( .A(\ab[29][13] ), .B(\CARRYB[28][13] ), .CI(\SUMB[28][14] ), 
        .CO(\CARRYB[29][13] ), .S(\SUMB[29][13] ) );
  FA_X1 S2_29_14 ( .A(\ab[29][14] ), .B(\CARRYB[28][14] ), .CI(\SUMB[28][15] ), 
        .CO(\CARRYB[29][14] ), .S(\SUMB[29][14] ) );
  FA_X1 S2_29_15 ( .A(\ab[29][15] ), .B(\CARRYB[28][15] ), .CI(\SUMB[28][16] ), 
        .CO(\CARRYB[29][15] ), .S(\SUMB[29][15] ) );
  FA_X1 S2_29_16 ( .A(\ab[29][16] ), .B(\CARRYB[28][16] ), .CI(\SUMB[28][17] ), 
        .CO(\CARRYB[29][16] ), .S(\SUMB[29][16] ) );
  FA_X1 S2_29_17 ( .A(\ab[29][17] ), .B(\CARRYB[28][17] ), .CI(\SUMB[28][18] ), 
        .CO(\CARRYB[29][17] ), .S(\SUMB[29][17] ) );
  FA_X1 S2_29_18 ( .A(\ab[29][18] ), .B(\CARRYB[28][18] ), .CI(\SUMB[28][19] ), 
        .CO(\CARRYB[29][18] ), .S(\SUMB[29][18] ) );
  FA_X1 S2_29_19 ( .A(\ab[29][19] ), .B(\CARRYB[28][19] ), .CI(\SUMB[28][20] ), 
        .CO(\CARRYB[29][19] ), .S(\SUMB[29][19] ) );
  FA_X1 S2_29_20 ( .A(\ab[29][20] ), .B(\CARRYB[28][20] ), .CI(\SUMB[28][21] ), 
        .CO(\CARRYB[29][20] ), .S(\SUMB[29][20] ) );
  FA_X1 S2_29_21 ( .A(\ab[29][21] ), .B(\CARRYB[28][21] ), .CI(\SUMB[28][22] ), 
        .CO(\CARRYB[29][21] ), .S(\SUMB[29][21] ) );
  FA_X1 S2_29_22 ( .A(\ab[29][22] ), .B(\CARRYB[28][22] ), .CI(\SUMB[28][23] ), 
        .CO(\CARRYB[29][22] ), .S(\SUMB[29][22] ) );
  FA_X1 S2_29_23 ( .A(\ab[29][23] ), .B(\CARRYB[28][23] ), .CI(\SUMB[28][24] ), 
        .CO(\CARRYB[29][23] ), .S(\SUMB[29][23] ) );
  FA_X1 S2_29_24 ( .A(\ab[29][24] ), .B(\CARRYB[28][24] ), .CI(\SUMB[28][25] ), 
        .CO(\CARRYB[29][24] ), .S(\SUMB[29][24] ) );
  FA_X1 S2_29_25 ( .A(\ab[29][25] ), .B(\CARRYB[28][25] ), .CI(\SUMB[28][26] ), 
        .CO(\CARRYB[29][25] ), .S(\SUMB[29][25] ) );
  FA_X1 S2_29_26 ( .A(\ab[29][26] ), .B(\CARRYB[28][26] ), .CI(\SUMB[28][27] ), 
        .CO(\CARRYB[29][26] ), .S(\SUMB[29][26] ) );
  FA_X1 S2_29_27 ( .A(\ab[29][27] ), .B(\CARRYB[28][27] ), .CI(\SUMB[28][28] ), 
        .CO(\CARRYB[29][27] ), .S(\SUMB[29][27] ) );
  FA_X1 S2_29_28 ( .A(\ab[29][28] ), .B(\CARRYB[28][28] ), .CI(\SUMB[28][29] ), 
        .CO(\CARRYB[29][28] ), .S(\SUMB[29][28] ) );
  FA_X1 S2_29_29 ( .A(\ab[29][29] ), .B(\CARRYB[28][29] ), .CI(\SUMB[28][30] ), 
        .CO(\CARRYB[29][29] ), .S(\SUMB[29][29] ) );
  FA_X1 S3_29_30 ( .A(\ab[29][30] ), .B(\CARRYB[28][30] ), .CI(\ab[28][31] ), 
        .CO(\CARRYB[29][30] ), .S(\SUMB[29][30] ) );
  FA_X1 S1_28_0 ( .A(\ab[28][0] ), .B(\CARRYB[27][0] ), .CI(\SUMB[27][1] ), 
        .CO(\CARRYB[28][0] ), .S(\A1[26] ) );
  FA_X1 S2_28_1 ( .A(\ab[28][1] ), .B(\CARRYB[27][1] ), .CI(\SUMB[27][2] ), 
        .CO(\CARRYB[28][1] ), .S(\SUMB[28][1] ) );
  FA_X1 S2_28_2 ( .A(\ab[28][2] ), .B(\CARRYB[27][2] ), .CI(\SUMB[27][3] ), 
        .CO(\CARRYB[28][2] ), .S(\SUMB[28][2] ) );
  FA_X1 S2_28_3 ( .A(\CARRYB[27][3] ), .B(\ab[28][3] ), .CI(\SUMB[27][4] ), 
        .CO(\CARRYB[28][3] ), .S(\SUMB[28][3] ) );
  FA_X1 S2_28_4 ( .A(\ab[28][4] ), .B(\CARRYB[27][4] ), .CI(\SUMB[27][5] ), 
        .CO(\CARRYB[28][4] ), .S(\SUMB[28][4] ) );
  FA_X1 S2_28_5 ( .A(\CARRYB[27][5] ), .B(\ab[28][5] ), .CI(\SUMB[27][6] ), 
        .CO(\CARRYB[28][5] ), .S(\SUMB[28][5] ) );
  FA_X1 S2_28_6 ( .A(\ab[28][6] ), .B(\CARRYB[27][6] ), .CI(\SUMB[27][7] ), 
        .CO(\CARRYB[28][6] ), .S(\SUMB[28][6] ) );
  FA_X1 S2_28_7 ( .A(\CARRYB[27][7] ), .B(\ab[28][7] ), .CI(\SUMB[27][8] ), 
        .CO(\CARRYB[28][7] ), .S(\SUMB[28][7] ) );
  FA_X1 S2_28_8 ( .A(\ab[28][8] ), .B(\CARRYB[27][8] ), .CI(\SUMB[27][9] ), 
        .CO(\CARRYB[28][8] ), .S(\SUMB[28][8] ) );
  FA_X1 S2_28_9 ( .A(\ab[28][9] ), .B(\CARRYB[27][9] ), .CI(\SUMB[27][10] ), 
        .CO(\CARRYB[28][9] ), .S(\SUMB[28][9] ) );
  FA_X1 S2_28_10 ( .A(\ab[28][10] ), .B(\CARRYB[27][10] ), .CI(\SUMB[27][11] ), 
        .CO(\CARRYB[28][10] ), .S(\SUMB[28][10] ) );
  FA_X1 S2_28_11 ( .A(\ab[28][11] ), .B(\CARRYB[27][11] ), .CI(\SUMB[27][12] ), 
        .CO(\CARRYB[28][11] ), .S(\SUMB[28][11] ) );
  FA_X1 S2_28_12 ( .A(\ab[28][12] ), .B(\CARRYB[27][12] ), .CI(\SUMB[27][13] ), 
        .CO(\CARRYB[28][12] ), .S(\SUMB[28][12] ) );
  FA_X1 S2_28_13 ( .A(\ab[28][13] ), .B(\CARRYB[27][13] ), .CI(\SUMB[27][14] ), 
        .CO(\CARRYB[28][13] ), .S(\SUMB[28][13] ) );
  FA_X1 S2_28_14 ( .A(\ab[28][14] ), .B(\CARRYB[27][14] ), .CI(\SUMB[27][15] ), 
        .CO(\CARRYB[28][14] ), .S(\SUMB[28][14] ) );
  FA_X1 S2_28_15 ( .A(\ab[28][15] ), .B(\CARRYB[27][15] ), .CI(\SUMB[27][16] ), 
        .CO(\CARRYB[28][15] ), .S(\SUMB[28][15] ) );
  FA_X1 S2_28_16 ( .A(\ab[28][16] ), .B(\CARRYB[27][16] ), .CI(\SUMB[27][17] ), 
        .CO(\CARRYB[28][16] ), .S(\SUMB[28][16] ) );
  FA_X1 S2_28_17 ( .A(\ab[28][17] ), .B(\CARRYB[27][17] ), .CI(\SUMB[27][18] ), 
        .CO(\CARRYB[28][17] ), .S(\SUMB[28][17] ) );
  FA_X1 S2_28_18 ( .A(\ab[28][18] ), .B(\CARRYB[27][18] ), .CI(\SUMB[27][19] ), 
        .CO(\CARRYB[28][18] ), .S(\SUMB[28][18] ) );
  FA_X1 S2_28_19 ( .A(\ab[28][19] ), .B(\CARRYB[27][19] ), .CI(\SUMB[27][20] ), 
        .CO(\CARRYB[28][19] ), .S(\SUMB[28][19] ) );
  FA_X1 S2_28_20 ( .A(\ab[28][20] ), .B(\CARRYB[27][20] ), .CI(\SUMB[27][21] ), 
        .CO(\CARRYB[28][20] ), .S(\SUMB[28][20] ) );
  FA_X1 S2_28_21 ( .A(\ab[28][21] ), .B(\CARRYB[27][21] ), .CI(\SUMB[27][22] ), 
        .CO(\CARRYB[28][21] ), .S(\SUMB[28][21] ) );
  FA_X1 S2_28_22 ( .A(\ab[28][22] ), .B(\CARRYB[27][22] ), .CI(\SUMB[27][23] ), 
        .CO(\CARRYB[28][22] ), .S(\SUMB[28][22] ) );
  FA_X1 S2_28_23 ( .A(\ab[28][23] ), .B(\CARRYB[27][23] ), .CI(\SUMB[27][24] ), 
        .CO(\CARRYB[28][23] ), .S(\SUMB[28][23] ) );
  FA_X1 S2_28_24 ( .A(\ab[28][24] ), .B(\CARRYB[27][24] ), .CI(\SUMB[27][25] ), 
        .CO(\CARRYB[28][24] ), .S(\SUMB[28][24] ) );
  FA_X1 S2_28_25 ( .A(\ab[28][25] ), .B(\CARRYB[27][25] ), .CI(\SUMB[27][26] ), 
        .CO(\CARRYB[28][25] ), .S(\SUMB[28][25] ) );
  FA_X1 S2_28_26 ( .A(\ab[28][26] ), .B(\CARRYB[27][26] ), .CI(\SUMB[27][27] ), 
        .CO(\CARRYB[28][26] ), .S(\SUMB[28][26] ) );
  FA_X1 S2_28_27 ( .A(\ab[28][27] ), .B(\CARRYB[27][27] ), .CI(\SUMB[27][28] ), 
        .CO(\CARRYB[28][27] ), .S(\SUMB[28][27] ) );
  FA_X1 S2_28_28 ( .A(\ab[28][28] ), .B(\CARRYB[27][28] ), .CI(\SUMB[27][29] ), 
        .CO(\CARRYB[28][28] ), .S(\SUMB[28][28] ) );
  FA_X1 S2_28_29 ( .A(\ab[28][29] ), .B(\CARRYB[27][29] ), .CI(\SUMB[27][30] ), 
        .CO(\CARRYB[28][29] ), .S(\SUMB[28][29] ) );
  FA_X1 S3_28_30 ( .A(\ab[28][30] ), .B(\CARRYB[27][30] ), .CI(\ab[27][31] ), 
        .CO(\CARRYB[28][30] ), .S(\SUMB[28][30] ) );
  FA_X1 S1_27_0 ( .A(\ab[27][0] ), .B(\CARRYB[26][0] ), .CI(\SUMB[26][1] ), 
        .CO(\CARRYB[27][0] ), .S(\A1[25] ) );
  FA_X1 S2_27_1 ( .A(\ab[27][1] ), .B(\CARRYB[26][1] ), .CI(\SUMB[26][2] ), 
        .CO(\CARRYB[27][1] ), .S(\SUMB[27][1] ) );
  FA_X1 S2_27_2 ( .A(\ab[27][2] ), .B(\CARRYB[26][2] ), .CI(\SUMB[26][3] ), 
        .CO(\CARRYB[27][2] ), .S(\SUMB[27][2] ) );
  FA_X1 S2_27_3 ( .A(\ab[27][3] ), .B(\CARRYB[26][3] ), .CI(\SUMB[26][4] ), 
        .CO(\CARRYB[27][3] ), .S(\SUMB[27][3] ) );
  FA_X1 S2_27_4 ( .A(\ab[27][4] ), .B(\CARRYB[26][4] ), .CI(\SUMB[26][5] ), 
        .CO(\CARRYB[27][4] ), .S(\SUMB[27][4] ) );
  FA_X1 S2_27_5 ( .A(\ab[27][5] ), .B(\CARRYB[26][5] ), .CI(\SUMB[26][6] ), 
        .CO(\CARRYB[27][5] ), .S(\SUMB[27][5] ) );
  FA_X1 S2_27_6 ( .A(\CARRYB[26][6] ), .B(\ab[27][6] ), .CI(\SUMB[26][7] ), 
        .CO(\CARRYB[27][6] ), .S(\SUMB[27][6] ) );
  FA_X1 S2_27_7 ( .A(\CARRYB[26][7] ), .B(\ab[27][7] ), .CI(\SUMB[26][8] ), 
        .CO(\CARRYB[27][7] ), .S(\SUMB[27][7] ) );
  FA_X1 S2_27_8 ( .A(\ab[27][8] ), .B(\CARRYB[26][8] ), .CI(\SUMB[26][9] ), 
        .CO(\CARRYB[27][8] ), .S(\SUMB[27][8] ) );
  FA_X1 S2_27_9 ( .A(\ab[27][9] ), .B(\CARRYB[26][9] ), .CI(\SUMB[26][10] ), 
        .CO(\CARRYB[27][9] ), .S(\SUMB[27][9] ) );
  FA_X1 S2_27_10 ( .A(\ab[27][10] ), .B(\CARRYB[26][10] ), .CI(\SUMB[26][11] ), 
        .CO(\CARRYB[27][10] ), .S(\SUMB[27][10] ) );
  FA_X1 S2_27_11 ( .A(\ab[27][11] ), .B(\CARRYB[26][11] ), .CI(\SUMB[26][12] ), 
        .CO(\CARRYB[27][11] ), .S(\SUMB[27][11] ) );
  FA_X1 S2_27_12 ( .A(\ab[27][12] ), .B(\CARRYB[26][12] ), .CI(\SUMB[26][13] ), 
        .CO(\CARRYB[27][12] ), .S(\SUMB[27][12] ) );
  FA_X1 S2_27_13 ( .A(\ab[27][13] ), .B(\CARRYB[26][13] ), .CI(\SUMB[26][14] ), 
        .CO(\CARRYB[27][13] ), .S(\SUMB[27][13] ) );
  FA_X1 S2_27_14 ( .A(\ab[27][14] ), .B(\CARRYB[26][14] ), .CI(\SUMB[26][15] ), 
        .CO(\CARRYB[27][14] ), .S(\SUMB[27][14] ) );
  FA_X1 S2_27_15 ( .A(\ab[27][15] ), .B(\CARRYB[26][15] ), .CI(\SUMB[26][16] ), 
        .CO(\CARRYB[27][15] ), .S(\SUMB[27][15] ) );
  FA_X1 S2_27_16 ( .A(\ab[27][16] ), .B(\CARRYB[26][16] ), .CI(\SUMB[26][17] ), 
        .CO(\CARRYB[27][16] ), .S(\SUMB[27][16] ) );
  FA_X1 S2_27_17 ( .A(\ab[27][17] ), .B(\CARRYB[26][17] ), .CI(\SUMB[26][18] ), 
        .CO(\CARRYB[27][17] ), .S(\SUMB[27][17] ) );
  FA_X1 S2_27_18 ( .A(\ab[27][18] ), .B(\CARRYB[26][18] ), .CI(\SUMB[26][19] ), 
        .CO(\CARRYB[27][18] ), .S(\SUMB[27][18] ) );
  FA_X1 S2_27_19 ( .A(\ab[27][19] ), .B(\CARRYB[26][19] ), .CI(\SUMB[26][20] ), 
        .CO(\CARRYB[27][19] ), .S(\SUMB[27][19] ) );
  FA_X1 S2_27_20 ( .A(\ab[27][20] ), .B(\CARRYB[26][20] ), .CI(\SUMB[26][21] ), 
        .CO(\CARRYB[27][20] ), .S(\SUMB[27][20] ) );
  FA_X1 S2_27_21 ( .A(\ab[27][21] ), .B(\CARRYB[26][21] ), .CI(\SUMB[26][22] ), 
        .CO(\CARRYB[27][21] ), .S(\SUMB[27][21] ) );
  FA_X1 S2_27_22 ( .A(\ab[27][22] ), .B(\CARRYB[26][22] ), .CI(\SUMB[26][23] ), 
        .CO(\CARRYB[27][22] ), .S(\SUMB[27][22] ) );
  FA_X1 S2_27_23 ( .A(\ab[27][23] ), .B(\CARRYB[26][23] ), .CI(\SUMB[26][24] ), 
        .CO(\CARRYB[27][23] ), .S(\SUMB[27][23] ) );
  FA_X1 S2_27_24 ( .A(\ab[27][24] ), .B(\CARRYB[26][24] ), .CI(\SUMB[26][25] ), 
        .CO(\CARRYB[27][24] ), .S(\SUMB[27][24] ) );
  FA_X1 S2_27_25 ( .A(\ab[27][25] ), .B(\CARRYB[26][25] ), .CI(\SUMB[26][26] ), 
        .CO(\CARRYB[27][25] ), .S(\SUMB[27][25] ) );
  FA_X1 S2_27_26 ( .A(\ab[27][26] ), .B(\CARRYB[26][26] ), .CI(\SUMB[26][27] ), 
        .CO(\CARRYB[27][26] ), .S(\SUMB[27][26] ) );
  FA_X1 S2_27_27 ( .A(\ab[27][27] ), .B(\CARRYB[26][27] ), .CI(\SUMB[26][28] ), 
        .CO(\CARRYB[27][27] ), .S(\SUMB[27][27] ) );
  FA_X1 S2_27_28 ( .A(\ab[27][28] ), .B(\CARRYB[26][28] ), .CI(\SUMB[26][29] ), 
        .CO(\CARRYB[27][28] ), .S(\SUMB[27][28] ) );
  FA_X1 S2_27_29 ( .A(\ab[27][29] ), .B(\CARRYB[26][29] ), .CI(\SUMB[26][30] ), 
        .CO(\CARRYB[27][29] ), .S(\SUMB[27][29] ) );
  FA_X1 S3_27_30 ( .A(\ab[27][30] ), .B(\CARRYB[26][30] ), .CI(\ab[26][31] ), 
        .CO(\CARRYB[27][30] ), .S(\SUMB[27][30] ) );
  FA_X1 S1_26_0 ( .A(\ab[26][0] ), .B(\CARRYB[25][0] ), .CI(\SUMB[25][1] ), 
        .CO(\CARRYB[26][0] ), .S(\A1[24] ) );
  FA_X1 S2_26_1 ( .A(\ab[26][1] ), .B(\CARRYB[25][1] ), .CI(\SUMB[25][2] ), 
        .CO(\CARRYB[26][1] ), .S(\SUMB[26][1] ) );
  FA_X1 S2_26_2 ( .A(\ab[26][2] ), .B(\CARRYB[25][2] ), .CI(\SUMB[25][3] ), 
        .CO(\CARRYB[26][2] ), .S(\SUMB[26][2] ) );
  FA_X1 S2_26_3 ( .A(\ab[26][3] ), .B(\CARRYB[25][3] ), .CI(\SUMB[25][4] ), 
        .CO(\CARRYB[26][3] ), .S(\SUMB[26][3] ) );
  FA_X1 S2_26_4 ( .A(\ab[26][4] ), .B(\CARRYB[25][4] ), .CI(\SUMB[25][5] ), 
        .CO(\CARRYB[26][4] ), .S(\SUMB[26][4] ) );
  FA_X1 S2_26_5 ( .A(\CARRYB[25][5] ), .B(\ab[26][5] ), .CI(\SUMB[25][6] ), 
        .CO(\CARRYB[26][5] ), .S(\SUMB[26][5] ) );
  FA_X1 S2_26_6 ( .A(\ab[26][6] ), .B(\CARRYB[25][6] ), .CI(\SUMB[25][7] ), 
        .CO(\CARRYB[26][6] ), .S(\SUMB[26][6] ) );
  FA_X1 S2_26_7 ( .A(\ab[26][7] ), .B(\CARRYB[25][7] ), .CI(\SUMB[25][8] ), 
        .CO(\CARRYB[26][7] ), .S(\SUMB[26][7] ) );
  FA_X1 S2_26_8 ( .A(\CARRYB[25][8] ), .B(\ab[26][8] ), .CI(\SUMB[25][9] ), 
        .CO(\CARRYB[26][8] ), .S(\SUMB[26][8] ) );
  FA_X1 S2_26_9 ( .A(\CARRYB[25][9] ), .B(\ab[26][9] ), .CI(\SUMB[25][10] ), 
        .CO(\CARRYB[26][9] ), .S(\SUMB[26][9] ) );
  FA_X1 S2_26_10 ( .A(\ab[26][10] ), .B(\CARRYB[25][10] ), .CI(\SUMB[25][11] ), 
        .CO(\CARRYB[26][10] ), .S(\SUMB[26][10] ) );
  FA_X1 S2_26_11 ( .A(\ab[26][11] ), .B(\CARRYB[25][11] ), .CI(\SUMB[25][12] ), 
        .CO(\CARRYB[26][11] ), .S(\SUMB[26][11] ) );
  FA_X1 S2_26_12 ( .A(\ab[26][12] ), .B(\CARRYB[25][12] ), .CI(\SUMB[25][13] ), 
        .CO(\CARRYB[26][12] ), .S(\SUMB[26][12] ) );
  FA_X1 S2_26_13 ( .A(\ab[26][13] ), .B(\CARRYB[25][13] ), .CI(\SUMB[25][14] ), 
        .CO(\CARRYB[26][13] ), .S(\SUMB[26][13] ) );
  FA_X1 S2_26_14 ( .A(\ab[26][14] ), .B(\CARRYB[25][14] ), .CI(\SUMB[25][15] ), 
        .CO(\CARRYB[26][14] ), .S(\SUMB[26][14] ) );
  FA_X1 S2_26_15 ( .A(\ab[26][15] ), .B(\CARRYB[25][15] ), .CI(\SUMB[25][16] ), 
        .CO(\CARRYB[26][15] ), .S(\SUMB[26][15] ) );
  FA_X1 S2_26_16 ( .A(\ab[26][16] ), .B(\CARRYB[25][16] ), .CI(\SUMB[25][17] ), 
        .CO(\CARRYB[26][16] ), .S(\SUMB[26][16] ) );
  FA_X1 S2_26_17 ( .A(\ab[26][17] ), .B(\CARRYB[25][17] ), .CI(\SUMB[25][18] ), 
        .CO(\CARRYB[26][17] ), .S(\SUMB[26][17] ) );
  FA_X1 S2_26_18 ( .A(\ab[26][18] ), .B(\CARRYB[25][18] ), .CI(\SUMB[25][19] ), 
        .CO(\CARRYB[26][18] ), .S(\SUMB[26][18] ) );
  FA_X1 S2_26_19 ( .A(\ab[26][19] ), .B(\CARRYB[25][19] ), .CI(\SUMB[25][20] ), 
        .CO(\CARRYB[26][19] ), .S(\SUMB[26][19] ) );
  FA_X1 S2_26_20 ( .A(\ab[26][20] ), .B(\CARRYB[25][20] ), .CI(\SUMB[25][21] ), 
        .CO(\CARRYB[26][20] ), .S(\SUMB[26][20] ) );
  FA_X1 S2_26_21 ( .A(\ab[26][21] ), .B(\CARRYB[25][21] ), .CI(\SUMB[25][22] ), 
        .CO(\CARRYB[26][21] ), .S(\SUMB[26][21] ) );
  FA_X1 S2_26_22 ( .A(\ab[26][22] ), .B(\CARRYB[25][22] ), .CI(\SUMB[25][23] ), 
        .CO(\CARRYB[26][22] ), .S(\SUMB[26][22] ) );
  FA_X1 S2_26_23 ( .A(\ab[26][23] ), .B(\CARRYB[25][23] ), .CI(\SUMB[25][24] ), 
        .CO(\CARRYB[26][23] ), .S(\SUMB[26][23] ) );
  FA_X1 S2_26_24 ( .A(\ab[26][24] ), .B(\CARRYB[25][24] ), .CI(\SUMB[25][25] ), 
        .CO(\CARRYB[26][24] ), .S(\SUMB[26][24] ) );
  FA_X1 S2_26_25 ( .A(\ab[26][25] ), .B(\CARRYB[25][25] ), .CI(\SUMB[25][26] ), 
        .CO(\CARRYB[26][25] ), .S(\SUMB[26][25] ) );
  FA_X1 S2_26_26 ( .A(\ab[26][26] ), .B(\CARRYB[25][26] ), .CI(\SUMB[25][27] ), 
        .CO(\CARRYB[26][26] ), .S(\SUMB[26][26] ) );
  FA_X1 S2_26_27 ( .A(\ab[26][27] ), .B(\CARRYB[25][27] ), .CI(\SUMB[25][28] ), 
        .CO(\CARRYB[26][27] ), .S(\SUMB[26][27] ) );
  FA_X1 S2_26_28 ( .A(\ab[26][28] ), .B(\CARRYB[25][28] ), .CI(\SUMB[25][29] ), 
        .CO(\CARRYB[26][28] ), .S(\SUMB[26][28] ) );
  FA_X1 S2_26_29 ( .A(\ab[26][29] ), .B(\CARRYB[25][29] ), .CI(\SUMB[25][30] ), 
        .CO(\CARRYB[26][29] ), .S(\SUMB[26][29] ) );
  FA_X1 S3_26_30 ( .A(\ab[26][30] ), .B(\CARRYB[25][30] ), .CI(\ab[25][31] ), 
        .CO(\CARRYB[26][30] ), .S(\SUMB[26][30] ) );
  FA_X1 S1_25_0 ( .A(\ab[25][0] ), .B(\CARRYB[24][0] ), .CI(\SUMB[24][1] ), 
        .CO(\CARRYB[25][0] ), .S(\A1[23] ) );
  FA_X1 S2_25_1 ( .A(\ab[25][1] ), .B(\CARRYB[24][1] ), .CI(\SUMB[24][2] ), 
        .CO(\CARRYB[25][1] ), .S(\SUMB[25][1] ) );
  FA_X1 S2_25_2 ( .A(\ab[25][2] ), .B(\CARRYB[24][2] ), .CI(\SUMB[24][3] ), 
        .CO(\CARRYB[25][2] ), .S(\SUMB[25][2] ) );
  FA_X1 S2_25_3 ( .A(\ab[25][3] ), .B(\CARRYB[24][3] ), .CI(\SUMB[24][4] ), 
        .CO(\CARRYB[25][3] ), .S(\SUMB[25][3] ) );
  FA_X1 S2_25_4 ( .A(\ab[25][4] ), .B(\CARRYB[24][4] ), .CI(\SUMB[24][5] ), 
        .CO(\CARRYB[25][4] ), .S(\SUMB[25][4] ) );
  FA_X1 S2_25_5 ( .A(\ab[25][5] ), .B(\CARRYB[24][5] ), .CI(\SUMB[24][6] ), 
        .CO(\CARRYB[25][5] ), .S(\SUMB[25][5] ) );
  FA_X1 S2_25_6 ( .A(\ab[25][6] ), .B(\CARRYB[24][6] ), .CI(\SUMB[24][7] ), 
        .CO(\CARRYB[25][6] ), .S(\SUMB[25][6] ) );
  FA_X1 S2_25_7 ( .A(\ab[25][7] ), .B(\CARRYB[24][7] ), .CI(\SUMB[24][8] ), 
        .CO(\CARRYB[25][7] ), .S(\SUMB[25][7] ) );
  FA_X1 S2_25_8 ( .A(\CARRYB[24][8] ), .B(\ab[25][8] ), .CI(\SUMB[24][9] ), 
        .CO(\CARRYB[25][8] ), .S(\SUMB[25][8] ) );
  FA_X1 S2_25_9 ( .A(\CARRYB[24][9] ), .B(\ab[25][9] ), .CI(\SUMB[24][10] ), 
        .CO(\CARRYB[25][9] ), .S(\SUMB[25][9] ) );
  FA_X1 S2_25_10 ( .A(\ab[25][10] ), .B(\CARRYB[24][10] ), .CI(\SUMB[24][11] ), 
        .CO(\CARRYB[25][10] ), .S(\SUMB[25][10] ) );
  FA_X1 S2_25_11 ( .A(\ab[25][11] ), .B(\CARRYB[24][11] ), .CI(\SUMB[24][12] ), 
        .CO(\CARRYB[25][11] ), .S(\SUMB[25][11] ) );
  FA_X1 S2_25_12 ( .A(\ab[25][12] ), .B(\CARRYB[24][12] ), .CI(\SUMB[24][13] ), 
        .CO(\CARRYB[25][12] ), .S(\SUMB[25][12] ) );
  FA_X1 S2_25_13 ( .A(\ab[25][13] ), .B(\CARRYB[24][13] ), .CI(\SUMB[24][14] ), 
        .CO(\CARRYB[25][13] ), .S(\SUMB[25][13] ) );
  FA_X1 S2_25_14 ( .A(\ab[25][14] ), .B(\CARRYB[24][14] ), .CI(\SUMB[24][15] ), 
        .CO(\CARRYB[25][14] ), .S(\SUMB[25][14] ) );
  FA_X1 S2_25_15 ( .A(\ab[25][15] ), .B(\CARRYB[24][15] ), .CI(\SUMB[24][16] ), 
        .CO(\CARRYB[25][15] ), .S(\SUMB[25][15] ) );
  FA_X1 S2_25_16 ( .A(\ab[25][16] ), .B(\CARRYB[24][16] ), .CI(\SUMB[24][17] ), 
        .CO(\CARRYB[25][16] ), .S(\SUMB[25][16] ) );
  FA_X1 S2_25_17 ( .A(\ab[25][17] ), .B(\CARRYB[24][17] ), .CI(\SUMB[24][18] ), 
        .CO(\CARRYB[25][17] ), .S(\SUMB[25][17] ) );
  FA_X1 S2_25_18 ( .A(\ab[25][18] ), .B(\CARRYB[24][18] ), .CI(\SUMB[24][19] ), 
        .CO(\CARRYB[25][18] ), .S(\SUMB[25][18] ) );
  FA_X1 S2_25_19 ( .A(\ab[25][19] ), .B(\CARRYB[24][19] ), .CI(\SUMB[24][20] ), 
        .CO(\CARRYB[25][19] ), .S(\SUMB[25][19] ) );
  FA_X1 S2_25_20 ( .A(\ab[25][20] ), .B(\CARRYB[24][20] ), .CI(\SUMB[24][21] ), 
        .CO(\CARRYB[25][20] ), .S(\SUMB[25][20] ) );
  FA_X1 S2_25_21 ( .A(\ab[25][21] ), .B(\CARRYB[24][21] ), .CI(\SUMB[24][22] ), 
        .CO(\CARRYB[25][21] ), .S(\SUMB[25][21] ) );
  FA_X1 S2_25_22 ( .A(\ab[25][22] ), .B(\CARRYB[24][22] ), .CI(\SUMB[24][23] ), 
        .CO(\CARRYB[25][22] ), .S(\SUMB[25][22] ) );
  FA_X1 S2_25_23 ( .A(\ab[25][23] ), .B(\CARRYB[24][23] ), .CI(\SUMB[24][24] ), 
        .CO(\CARRYB[25][23] ), .S(\SUMB[25][23] ) );
  FA_X1 S2_25_24 ( .A(\ab[25][24] ), .B(\CARRYB[24][24] ), .CI(\SUMB[24][25] ), 
        .CO(\CARRYB[25][24] ), .S(\SUMB[25][24] ) );
  FA_X1 S2_25_25 ( .A(\ab[25][25] ), .B(\CARRYB[24][25] ), .CI(\SUMB[24][26] ), 
        .CO(\CARRYB[25][25] ), .S(\SUMB[25][25] ) );
  FA_X1 S2_25_26 ( .A(\ab[25][26] ), .B(\CARRYB[24][26] ), .CI(\SUMB[24][27] ), 
        .CO(\CARRYB[25][26] ), .S(\SUMB[25][26] ) );
  FA_X1 S2_25_27 ( .A(\ab[25][27] ), .B(\CARRYB[24][27] ), .CI(\SUMB[24][28] ), 
        .CO(\CARRYB[25][27] ), .S(\SUMB[25][27] ) );
  FA_X1 S2_25_28 ( .A(\ab[25][28] ), .B(\CARRYB[24][28] ), .CI(\SUMB[24][29] ), 
        .CO(\CARRYB[25][28] ), .S(\SUMB[25][28] ) );
  FA_X1 S2_25_29 ( .A(\ab[25][29] ), .B(\CARRYB[24][29] ), .CI(\SUMB[24][30] ), 
        .CO(\CARRYB[25][29] ), .S(\SUMB[25][29] ) );
  FA_X1 S3_25_30 ( .A(\ab[25][30] ), .B(\CARRYB[24][30] ), .CI(\ab[24][31] ), 
        .CO(\CARRYB[25][30] ), .S(\SUMB[25][30] ) );
  FA_X1 S1_24_0 ( .A(\ab[24][0] ), .B(\CARRYB[23][0] ), .CI(\SUMB[23][1] ), 
        .CO(\CARRYB[24][0] ), .S(\A1[22] ) );
  FA_X1 S2_24_1 ( .A(\ab[24][1] ), .B(\CARRYB[23][1] ), .CI(\SUMB[23][2] ), 
        .CO(\CARRYB[24][1] ), .S(\SUMB[24][1] ) );
  FA_X1 S2_24_2 ( .A(\ab[24][2] ), .B(\CARRYB[23][2] ), .CI(\SUMB[23][3] ), 
        .CO(\CARRYB[24][2] ), .S(\SUMB[24][2] ) );
  FA_X1 S2_24_3 ( .A(\ab[24][3] ), .B(\CARRYB[23][3] ), .CI(\SUMB[23][4] ), 
        .CO(\CARRYB[24][3] ), .S(\SUMB[24][3] ) );
  FA_X1 S2_24_4 ( .A(\ab[24][4] ), .B(\CARRYB[23][4] ), .CI(\SUMB[23][5] ), 
        .CO(\CARRYB[24][4] ), .S(\SUMB[24][4] ) );
  FA_X1 S2_24_5 ( .A(\ab[24][5] ), .B(\CARRYB[23][5] ), .CI(\SUMB[23][6] ), 
        .CO(\CARRYB[24][5] ), .S(\SUMB[24][5] ) );
  FA_X1 S2_24_6 ( .A(\ab[24][6] ), .B(\CARRYB[23][6] ), .CI(\SUMB[23][7] ), 
        .CO(\CARRYB[24][6] ), .S(\SUMB[24][6] ) );
  FA_X1 S2_24_7 ( .A(\ab[24][7] ), .B(\CARRYB[23][7] ), .CI(\SUMB[23][8] ), 
        .CO(\CARRYB[24][7] ), .S(\SUMB[24][7] ) );
  FA_X1 S2_24_8 ( .A(\ab[24][8] ), .B(\CARRYB[23][8] ), .CI(\SUMB[23][9] ), 
        .CO(\CARRYB[24][8] ), .S(\SUMB[24][8] ) );
  FA_X1 S2_24_9 ( .A(\ab[24][9] ), .B(\CARRYB[23][9] ), .CI(\SUMB[23][10] ), 
        .CO(\CARRYB[24][9] ), .S(\SUMB[24][9] ) );
  FA_X1 S2_24_10 ( .A(\ab[24][10] ), .B(\CARRYB[23][10] ), .CI(\SUMB[23][11] ), 
        .CO(\CARRYB[24][10] ), .S(\SUMB[24][10] ) );
  FA_X1 S2_24_11 ( .A(\CARRYB[23][11] ), .B(\ab[24][11] ), .CI(\SUMB[23][12] ), 
        .CO(\CARRYB[24][11] ), .S(\SUMB[24][11] ) );
  FA_X1 S2_24_12 ( .A(\ab[24][12] ), .B(\CARRYB[23][12] ), .CI(\SUMB[23][13] ), 
        .CO(\CARRYB[24][12] ), .S(\SUMB[24][12] ) );
  FA_X1 S2_24_13 ( .A(\ab[24][13] ), .B(\CARRYB[23][13] ), .CI(\SUMB[23][14] ), 
        .CO(\CARRYB[24][13] ), .S(\SUMB[24][13] ) );
  FA_X1 S2_24_14 ( .A(\ab[24][14] ), .B(\CARRYB[23][14] ), .CI(\SUMB[23][15] ), 
        .CO(\CARRYB[24][14] ), .S(\SUMB[24][14] ) );
  FA_X1 S2_24_15 ( .A(\ab[24][15] ), .B(\CARRYB[23][15] ), .CI(\SUMB[23][16] ), 
        .CO(\CARRYB[24][15] ), .S(\SUMB[24][15] ) );
  FA_X1 S2_24_16 ( .A(\ab[24][16] ), .B(\CARRYB[23][16] ), .CI(\SUMB[23][17] ), 
        .CO(\CARRYB[24][16] ), .S(\SUMB[24][16] ) );
  FA_X1 S2_24_17 ( .A(\ab[24][17] ), .B(\CARRYB[23][17] ), .CI(\SUMB[23][18] ), 
        .CO(\CARRYB[24][17] ), .S(\SUMB[24][17] ) );
  FA_X1 S2_24_18 ( .A(\ab[24][18] ), .B(\CARRYB[23][18] ), .CI(\SUMB[23][19] ), 
        .CO(\CARRYB[24][18] ), .S(\SUMB[24][18] ) );
  FA_X1 S2_24_19 ( .A(\ab[24][19] ), .B(\CARRYB[23][19] ), .CI(\SUMB[23][20] ), 
        .CO(\CARRYB[24][19] ), .S(\SUMB[24][19] ) );
  FA_X1 S2_24_20 ( .A(\ab[24][20] ), .B(\CARRYB[23][20] ), .CI(\SUMB[23][21] ), 
        .CO(\CARRYB[24][20] ), .S(\SUMB[24][20] ) );
  FA_X1 S2_24_21 ( .A(\ab[24][21] ), .B(\CARRYB[23][21] ), .CI(\SUMB[23][22] ), 
        .CO(\CARRYB[24][21] ), .S(\SUMB[24][21] ) );
  FA_X1 S2_24_22 ( .A(\ab[24][22] ), .B(\CARRYB[23][22] ), .CI(\SUMB[23][23] ), 
        .CO(\CARRYB[24][22] ), .S(\SUMB[24][22] ) );
  FA_X1 S2_24_23 ( .A(\ab[24][23] ), .B(\CARRYB[23][23] ), .CI(\SUMB[23][24] ), 
        .CO(\CARRYB[24][23] ), .S(\SUMB[24][23] ) );
  FA_X1 S2_24_24 ( .A(\ab[24][24] ), .B(\CARRYB[23][24] ), .CI(\SUMB[23][25] ), 
        .CO(\CARRYB[24][24] ), .S(\SUMB[24][24] ) );
  FA_X1 S2_24_25 ( .A(\ab[24][25] ), .B(\CARRYB[23][25] ), .CI(\SUMB[23][26] ), 
        .CO(\CARRYB[24][25] ), .S(\SUMB[24][25] ) );
  FA_X1 S2_24_26 ( .A(\ab[24][26] ), .B(\CARRYB[23][26] ), .CI(\SUMB[23][27] ), 
        .CO(\CARRYB[24][26] ), .S(\SUMB[24][26] ) );
  FA_X1 S2_24_27 ( .A(\ab[24][27] ), .B(\CARRYB[23][27] ), .CI(\SUMB[23][28] ), 
        .CO(\CARRYB[24][27] ), .S(\SUMB[24][27] ) );
  FA_X1 S2_24_28 ( .A(\ab[24][28] ), .B(\CARRYB[23][28] ), .CI(\SUMB[23][29] ), 
        .CO(\CARRYB[24][28] ), .S(\SUMB[24][28] ) );
  FA_X1 S2_24_29 ( .A(\ab[24][29] ), .B(\CARRYB[23][29] ), .CI(\SUMB[23][30] ), 
        .CO(\CARRYB[24][29] ), .S(\SUMB[24][29] ) );
  FA_X1 S3_24_30 ( .A(\ab[24][30] ), .B(\CARRYB[23][30] ), .CI(\ab[23][31] ), 
        .CO(\CARRYB[24][30] ), .S(\SUMB[24][30] ) );
  FA_X1 S1_23_0 ( .A(\ab[23][0] ), .B(\CARRYB[22][0] ), .CI(\SUMB[22][1] ), 
        .CO(\CARRYB[23][0] ), .S(\A1[21] ) );
  FA_X1 S2_23_1 ( .A(\ab[23][1] ), .B(\CARRYB[22][1] ), .CI(\SUMB[22][2] ), 
        .CO(\CARRYB[23][1] ), .S(\SUMB[23][1] ) );
  FA_X1 S2_23_2 ( .A(\ab[23][2] ), .B(\CARRYB[22][2] ), .CI(\SUMB[22][3] ), 
        .CO(\CARRYB[23][2] ), .S(\SUMB[23][2] ) );
  FA_X1 S2_23_3 ( .A(\ab[23][3] ), .B(\CARRYB[22][3] ), .CI(\SUMB[22][4] ), 
        .CO(\CARRYB[23][3] ), .S(\SUMB[23][3] ) );
  FA_X1 S2_23_4 ( .A(\ab[23][4] ), .B(\CARRYB[22][4] ), .CI(\SUMB[22][5] ), 
        .CO(\CARRYB[23][4] ), .S(\SUMB[23][4] ) );
  FA_X1 S2_23_5 ( .A(\ab[23][5] ), .B(\CARRYB[22][5] ), .CI(\SUMB[22][6] ), 
        .CO(\CARRYB[23][5] ), .S(\SUMB[23][5] ) );
  FA_X1 S2_23_6 ( .A(\ab[23][6] ), .B(\CARRYB[22][6] ), .CI(\SUMB[22][7] ), 
        .CO(\CARRYB[23][6] ), .S(\SUMB[23][6] ) );
  FA_X1 S2_23_7 ( .A(\ab[23][7] ), .B(\CARRYB[22][7] ), .CI(\SUMB[22][8] ), 
        .CO(\CARRYB[23][7] ), .S(\SUMB[23][7] ) );
  FA_X1 S2_23_8 ( .A(\ab[23][8] ), .B(\CARRYB[22][8] ), .CI(\SUMB[22][9] ), 
        .CO(\CARRYB[23][8] ), .S(\SUMB[23][8] ) );
  FA_X1 S2_23_9 ( .A(\ab[23][9] ), .B(\CARRYB[22][9] ), .CI(\SUMB[22][10] ), 
        .CO(\CARRYB[23][9] ), .S(\SUMB[23][9] ) );
  FA_X1 S2_23_10 ( .A(\CARRYB[22][10] ), .B(\ab[23][10] ), .CI(\SUMB[22][11] ), 
        .CO(\CARRYB[23][10] ), .S(\SUMB[23][10] ) );
  FA_X1 S2_23_11 ( .A(\CARRYB[22][11] ), .B(\ab[23][11] ), .CI(\SUMB[22][12] ), 
        .CO(\CARRYB[23][11] ), .S(\SUMB[23][11] ) );
  FA_X1 S2_23_12 ( .A(\ab[23][12] ), .B(\CARRYB[22][12] ), .CI(\SUMB[22][13] ), 
        .CO(\CARRYB[23][12] ), .S(\SUMB[23][12] ) );
  FA_X1 S2_23_13 ( .A(\ab[23][13] ), .B(\CARRYB[22][13] ), .CI(\SUMB[22][14] ), 
        .CO(\CARRYB[23][13] ), .S(\SUMB[23][13] ) );
  FA_X1 S2_23_14 ( .A(\ab[23][14] ), .B(\CARRYB[22][14] ), .CI(\SUMB[22][15] ), 
        .CO(\CARRYB[23][14] ), .S(\SUMB[23][14] ) );
  FA_X1 S2_23_15 ( .A(\ab[23][15] ), .B(\CARRYB[22][15] ), .CI(\SUMB[22][16] ), 
        .CO(\CARRYB[23][15] ), .S(\SUMB[23][15] ) );
  FA_X1 S2_23_16 ( .A(\ab[23][16] ), .B(\CARRYB[22][16] ), .CI(\SUMB[22][17] ), 
        .CO(\CARRYB[23][16] ), .S(\SUMB[23][16] ) );
  FA_X1 S2_23_17 ( .A(\ab[23][17] ), .B(\CARRYB[22][17] ), .CI(\SUMB[22][18] ), 
        .CO(\CARRYB[23][17] ), .S(\SUMB[23][17] ) );
  FA_X1 S2_23_18 ( .A(\ab[23][18] ), .B(\CARRYB[22][18] ), .CI(\SUMB[22][19] ), 
        .CO(\CARRYB[23][18] ), .S(\SUMB[23][18] ) );
  FA_X1 S2_23_19 ( .A(\ab[23][19] ), .B(\CARRYB[22][19] ), .CI(\SUMB[22][20] ), 
        .CO(\CARRYB[23][19] ), .S(\SUMB[23][19] ) );
  FA_X1 S2_23_20 ( .A(\ab[23][20] ), .B(\CARRYB[22][20] ), .CI(\SUMB[22][21] ), 
        .CO(\CARRYB[23][20] ), .S(\SUMB[23][20] ) );
  FA_X1 S2_23_21 ( .A(\ab[23][21] ), .B(\CARRYB[22][21] ), .CI(\SUMB[22][22] ), 
        .CO(\CARRYB[23][21] ), .S(\SUMB[23][21] ) );
  FA_X1 S2_23_22 ( .A(\ab[23][22] ), .B(\CARRYB[22][22] ), .CI(\SUMB[22][23] ), 
        .CO(\CARRYB[23][22] ), .S(\SUMB[23][22] ) );
  FA_X1 S2_23_23 ( .A(\ab[23][23] ), .B(\CARRYB[22][23] ), .CI(\SUMB[22][24] ), 
        .CO(\CARRYB[23][23] ), .S(\SUMB[23][23] ) );
  FA_X1 S2_23_24 ( .A(\ab[23][24] ), .B(\CARRYB[22][24] ), .CI(\SUMB[22][25] ), 
        .CO(\CARRYB[23][24] ), .S(\SUMB[23][24] ) );
  FA_X1 S2_23_25 ( .A(\ab[23][25] ), .B(\CARRYB[22][25] ), .CI(\SUMB[22][26] ), 
        .CO(\CARRYB[23][25] ), .S(\SUMB[23][25] ) );
  FA_X1 S2_23_26 ( .A(\ab[23][26] ), .B(\CARRYB[22][26] ), .CI(\SUMB[22][27] ), 
        .CO(\CARRYB[23][26] ), .S(\SUMB[23][26] ) );
  FA_X1 S2_23_27 ( .A(\ab[23][27] ), .B(\CARRYB[22][27] ), .CI(\SUMB[22][28] ), 
        .CO(\CARRYB[23][27] ), .S(\SUMB[23][27] ) );
  FA_X1 S2_23_28 ( .A(\ab[23][28] ), .B(\CARRYB[22][28] ), .CI(\SUMB[22][29] ), 
        .CO(\CARRYB[23][28] ), .S(\SUMB[23][28] ) );
  FA_X1 S2_23_29 ( .A(\ab[23][29] ), .B(\CARRYB[22][29] ), .CI(\SUMB[22][30] ), 
        .CO(\CARRYB[23][29] ), .S(\SUMB[23][29] ) );
  FA_X1 S3_23_30 ( .A(\ab[23][30] ), .B(\CARRYB[22][30] ), .CI(\ab[22][31] ), 
        .CO(\CARRYB[23][30] ), .S(\SUMB[23][30] ) );
  FA_X1 S1_22_0 ( .A(\ab[22][0] ), .B(\CARRYB[21][0] ), .CI(\SUMB[21][1] ), 
        .CO(\CARRYB[22][0] ), .S(\A1[20] ) );
  FA_X1 S2_22_1 ( .A(\ab[22][1] ), .B(\CARRYB[21][1] ), .CI(\SUMB[21][2] ), 
        .CO(\CARRYB[22][1] ), .S(\SUMB[22][1] ) );
  FA_X1 S2_22_2 ( .A(\ab[22][2] ), .B(\CARRYB[21][2] ), .CI(\SUMB[21][3] ), 
        .CO(\CARRYB[22][2] ), .S(\SUMB[22][2] ) );
  FA_X1 S2_22_3 ( .A(\ab[22][3] ), .B(\CARRYB[21][3] ), .CI(\SUMB[21][4] ), 
        .CO(\CARRYB[22][3] ), .S(\SUMB[22][3] ) );
  FA_X1 S2_22_4 ( .A(\ab[22][4] ), .B(\CARRYB[21][4] ), .CI(\SUMB[21][5] ), 
        .CO(\CARRYB[22][4] ), .S(\SUMB[22][4] ) );
  FA_X1 S2_22_5 ( .A(\ab[22][5] ), .B(\CARRYB[21][5] ), .CI(\SUMB[21][6] ), 
        .CO(\CARRYB[22][5] ), .S(\SUMB[22][5] ) );
  FA_X1 S2_22_6 ( .A(\ab[22][6] ), .B(\CARRYB[21][6] ), .CI(\SUMB[21][7] ), 
        .CO(\CARRYB[22][6] ), .S(\SUMB[22][6] ) );
  FA_X1 S2_22_7 ( .A(\ab[22][7] ), .B(\CARRYB[21][7] ), .CI(\SUMB[21][8] ), 
        .CO(\CARRYB[22][7] ), .S(\SUMB[22][7] ) );
  FA_X1 S2_22_8 ( .A(\ab[22][8] ), .B(\CARRYB[21][8] ), .CI(\SUMB[21][9] ), 
        .CO(\CARRYB[22][8] ), .S(\SUMB[22][8] ) );
  FA_X1 S2_22_9 ( .A(\ab[22][9] ), .B(\CARRYB[21][9] ), .CI(\SUMB[21][10] ), 
        .CO(\CARRYB[22][9] ), .S(\SUMB[22][9] ) );
  FA_X1 S2_22_10 ( .A(\ab[22][10] ), .B(\CARRYB[21][10] ), .CI(\SUMB[21][11] ), 
        .CO(\CARRYB[22][10] ), .S(\SUMB[22][10] ) );
  FA_X1 S2_22_11 ( .A(\ab[22][11] ), .B(\CARRYB[21][11] ), .CI(\SUMB[21][12] ), 
        .CO(\CARRYB[22][11] ), .S(\SUMB[22][11] ) );
  FA_X1 S2_22_12 ( .A(\ab[22][12] ), .B(\CARRYB[21][12] ), .CI(\SUMB[21][13] ), 
        .CO(\CARRYB[22][12] ), .S(\SUMB[22][12] ) );
  FA_X1 S2_22_13 ( .A(\CARRYB[21][13] ), .B(\ab[22][13] ), .CI(\SUMB[21][14] ), 
        .CO(\CARRYB[22][13] ), .S(\SUMB[22][13] ) );
  FA_X1 S2_22_14 ( .A(\ab[22][14] ), .B(\CARRYB[21][14] ), .CI(\SUMB[21][15] ), 
        .CO(\CARRYB[22][14] ), .S(\SUMB[22][14] ) );
  FA_X1 S2_22_15 ( .A(\ab[22][15] ), .B(\CARRYB[21][15] ), .CI(\SUMB[21][16] ), 
        .CO(\CARRYB[22][15] ), .S(\SUMB[22][15] ) );
  FA_X1 S2_22_16 ( .A(\ab[22][16] ), .B(\CARRYB[21][16] ), .CI(\SUMB[21][17] ), 
        .CO(\CARRYB[22][16] ), .S(\SUMB[22][16] ) );
  FA_X1 S2_22_17 ( .A(\ab[22][17] ), .B(\CARRYB[21][17] ), .CI(\SUMB[21][18] ), 
        .CO(\CARRYB[22][17] ), .S(\SUMB[22][17] ) );
  FA_X1 S2_22_18 ( .A(\ab[22][18] ), .B(\CARRYB[21][18] ), .CI(\SUMB[21][19] ), 
        .CO(\CARRYB[22][18] ), .S(\SUMB[22][18] ) );
  FA_X1 S2_22_19 ( .A(\ab[22][19] ), .B(\CARRYB[21][19] ), .CI(\SUMB[21][20] ), 
        .CO(\CARRYB[22][19] ), .S(\SUMB[22][19] ) );
  FA_X1 S2_22_20 ( .A(\ab[22][20] ), .B(\CARRYB[21][20] ), .CI(\SUMB[21][21] ), 
        .CO(\CARRYB[22][20] ), .S(\SUMB[22][20] ) );
  FA_X1 S2_22_21 ( .A(\ab[22][21] ), .B(\CARRYB[21][21] ), .CI(\SUMB[21][22] ), 
        .CO(\CARRYB[22][21] ), .S(\SUMB[22][21] ) );
  FA_X1 S2_22_22 ( .A(\ab[22][22] ), .B(\CARRYB[21][22] ), .CI(\SUMB[21][23] ), 
        .CO(\CARRYB[22][22] ), .S(\SUMB[22][22] ) );
  FA_X1 S2_22_23 ( .A(\ab[22][23] ), .B(\CARRYB[21][23] ), .CI(\SUMB[21][24] ), 
        .CO(\CARRYB[22][23] ), .S(\SUMB[22][23] ) );
  FA_X1 S2_22_24 ( .A(\ab[22][24] ), .B(\CARRYB[21][24] ), .CI(\SUMB[21][25] ), 
        .CO(\CARRYB[22][24] ), .S(\SUMB[22][24] ) );
  FA_X1 S2_22_25 ( .A(\ab[22][25] ), .B(\CARRYB[21][25] ), .CI(\SUMB[21][26] ), 
        .CO(\CARRYB[22][25] ), .S(\SUMB[22][25] ) );
  FA_X1 S2_22_26 ( .A(\ab[22][26] ), .B(\CARRYB[21][26] ), .CI(\SUMB[21][27] ), 
        .CO(\CARRYB[22][26] ), .S(\SUMB[22][26] ) );
  FA_X1 S2_22_27 ( .A(\ab[22][27] ), .B(\CARRYB[21][27] ), .CI(\SUMB[21][28] ), 
        .CO(\CARRYB[22][27] ), .S(\SUMB[22][27] ) );
  FA_X1 S2_22_28 ( .A(\ab[22][28] ), .B(\CARRYB[21][28] ), .CI(\SUMB[21][29] ), 
        .CO(\CARRYB[22][28] ), .S(\SUMB[22][28] ) );
  FA_X1 S2_22_29 ( .A(\ab[22][29] ), .B(\CARRYB[21][29] ), .CI(\SUMB[21][30] ), 
        .CO(\CARRYB[22][29] ), .S(\SUMB[22][29] ) );
  FA_X1 S3_22_30 ( .A(\ab[22][30] ), .B(\CARRYB[21][30] ), .CI(\ab[21][31] ), 
        .CO(\CARRYB[22][30] ), .S(\SUMB[22][30] ) );
  FA_X1 S1_21_0 ( .A(\ab[21][0] ), .B(\CARRYB[20][0] ), .CI(\SUMB[20][1] ), 
        .CO(\CARRYB[21][0] ), .S(\A1[19] ) );
  FA_X1 S2_21_1 ( .A(\ab[21][1] ), .B(\CARRYB[20][1] ), .CI(\SUMB[20][2] ), 
        .CO(\CARRYB[21][1] ), .S(\SUMB[21][1] ) );
  FA_X1 S2_21_2 ( .A(\ab[21][2] ), .B(\CARRYB[20][2] ), .CI(\SUMB[20][3] ), 
        .CO(\CARRYB[21][2] ), .S(\SUMB[21][2] ) );
  FA_X1 S2_21_3 ( .A(\ab[21][3] ), .B(\CARRYB[20][3] ), .CI(\SUMB[20][4] ), 
        .CO(\CARRYB[21][3] ), .S(\SUMB[21][3] ) );
  FA_X1 S2_21_4 ( .A(\ab[21][4] ), .B(\CARRYB[20][4] ), .CI(\SUMB[20][5] ), 
        .CO(\CARRYB[21][4] ), .S(\SUMB[21][4] ) );
  FA_X1 S2_21_5 ( .A(\ab[21][5] ), .B(\CARRYB[20][5] ), .CI(\SUMB[20][6] ), 
        .CO(\CARRYB[21][5] ), .S(\SUMB[21][5] ) );
  FA_X1 S2_21_6 ( .A(\ab[21][6] ), .B(\CARRYB[20][6] ), .CI(\SUMB[20][7] ), 
        .CO(\CARRYB[21][6] ), .S(\SUMB[21][6] ) );
  FA_X1 S2_21_7 ( .A(\ab[21][7] ), .B(\CARRYB[20][7] ), .CI(\SUMB[20][8] ), 
        .CO(\CARRYB[21][7] ), .S(\SUMB[21][7] ) );
  FA_X1 S2_21_8 ( .A(\ab[21][8] ), .B(\CARRYB[20][8] ), .CI(\SUMB[20][9] ), 
        .CO(\CARRYB[21][8] ), .S(\SUMB[21][8] ) );
  FA_X1 S2_21_9 ( .A(\CARRYB[20][9] ), .B(\ab[21][9] ), .CI(\SUMB[20][10] ), 
        .CO(\CARRYB[21][9] ), .S(\SUMB[21][9] ) );
  FA_X1 S2_21_10 ( .A(\ab[21][10] ), .B(\CARRYB[20][10] ), .CI(\SUMB[20][11] ), 
        .CO(\CARRYB[21][10] ), .S(\SUMB[21][10] ) );
  FA_X1 S2_21_11 ( .A(\ab[21][11] ), .B(\CARRYB[20][11] ), .CI(\SUMB[20][12] ), 
        .CO(\CARRYB[21][11] ), .S(\SUMB[21][11] ) );
  FA_X1 S2_21_12 ( .A(\ab[21][12] ), .B(\CARRYB[20][12] ), .CI(\SUMB[20][13] ), 
        .CO(\CARRYB[21][12] ), .S(\SUMB[21][12] ) );
  FA_X1 S2_21_13 ( .A(\CARRYB[20][13] ), .B(\ab[21][13] ), .CI(\SUMB[20][14] ), 
        .CO(\CARRYB[21][13] ), .S(\SUMB[21][13] ) );
  FA_X1 S2_21_14 ( .A(\ab[21][14] ), .B(\CARRYB[20][14] ), .CI(\SUMB[20][15] ), 
        .CO(\CARRYB[21][14] ), .S(\SUMB[21][14] ) );
  FA_X1 S2_21_15 ( .A(\ab[21][15] ), .B(\CARRYB[20][15] ), .CI(\SUMB[20][16] ), 
        .CO(\CARRYB[21][15] ), .S(\SUMB[21][15] ) );
  FA_X1 S2_21_16 ( .A(\ab[21][16] ), .B(\CARRYB[20][16] ), .CI(\SUMB[20][17] ), 
        .CO(\CARRYB[21][16] ), .S(\SUMB[21][16] ) );
  FA_X1 S2_21_17 ( .A(\ab[21][17] ), .B(\CARRYB[20][17] ), .CI(\SUMB[20][18] ), 
        .CO(\CARRYB[21][17] ), .S(\SUMB[21][17] ) );
  FA_X1 S2_21_18 ( .A(\ab[21][18] ), .B(\CARRYB[20][18] ), .CI(\SUMB[20][19] ), 
        .CO(\CARRYB[21][18] ), .S(\SUMB[21][18] ) );
  FA_X1 S2_21_19 ( .A(\ab[21][19] ), .B(\CARRYB[20][19] ), .CI(\SUMB[20][20] ), 
        .CO(\CARRYB[21][19] ), .S(\SUMB[21][19] ) );
  FA_X1 S2_21_20 ( .A(\ab[21][20] ), .B(\CARRYB[20][20] ), .CI(\SUMB[20][21] ), 
        .CO(\CARRYB[21][20] ), .S(\SUMB[21][20] ) );
  FA_X1 S2_21_21 ( .A(\ab[21][21] ), .B(\CARRYB[20][21] ), .CI(\SUMB[20][22] ), 
        .CO(\CARRYB[21][21] ), .S(\SUMB[21][21] ) );
  FA_X1 S2_21_22 ( .A(\ab[21][22] ), .B(\CARRYB[20][22] ), .CI(\SUMB[20][23] ), 
        .CO(\CARRYB[21][22] ), .S(\SUMB[21][22] ) );
  FA_X1 S2_21_23 ( .A(\ab[21][23] ), .B(\CARRYB[20][23] ), .CI(\SUMB[20][24] ), 
        .CO(\CARRYB[21][23] ), .S(\SUMB[21][23] ) );
  FA_X1 S2_21_24 ( .A(\ab[21][24] ), .B(\CARRYB[20][24] ), .CI(\SUMB[20][25] ), 
        .CO(\CARRYB[21][24] ), .S(\SUMB[21][24] ) );
  FA_X1 S2_21_25 ( .A(\ab[21][25] ), .B(\CARRYB[20][25] ), .CI(\SUMB[20][26] ), 
        .CO(\CARRYB[21][25] ), .S(\SUMB[21][25] ) );
  FA_X1 S2_21_26 ( .A(\ab[21][26] ), .B(\CARRYB[20][26] ), .CI(\SUMB[20][27] ), 
        .CO(\CARRYB[21][26] ), .S(\SUMB[21][26] ) );
  FA_X1 S2_21_27 ( .A(\ab[21][27] ), .B(\CARRYB[20][27] ), .CI(\SUMB[20][28] ), 
        .CO(\CARRYB[21][27] ), .S(\SUMB[21][27] ) );
  FA_X1 S2_21_28 ( .A(\ab[21][28] ), .B(\CARRYB[20][28] ), .CI(\SUMB[20][29] ), 
        .CO(\CARRYB[21][28] ), .S(\SUMB[21][28] ) );
  FA_X1 S2_21_29 ( .A(\ab[21][29] ), .B(\CARRYB[20][29] ), .CI(\SUMB[20][30] ), 
        .CO(\CARRYB[21][29] ), .S(\SUMB[21][29] ) );
  FA_X1 S3_21_30 ( .A(\ab[21][30] ), .B(\CARRYB[20][30] ), .CI(\ab[20][31] ), 
        .CO(\CARRYB[21][30] ), .S(\SUMB[21][30] ) );
  FA_X1 S1_20_0 ( .A(\ab[20][0] ), .B(\CARRYB[19][0] ), .CI(\SUMB[19][1] ), 
        .CO(\CARRYB[20][0] ), .S(\A1[18] ) );
  FA_X1 S2_20_1 ( .A(\ab[20][1] ), .B(\CARRYB[19][1] ), .CI(\SUMB[19][2] ), 
        .CO(\CARRYB[20][1] ), .S(\SUMB[20][1] ) );
  FA_X1 S2_20_2 ( .A(\ab[20][2] ), .B(\CARRYB[19][2] ), .CI(\SUMB[19][3] ), 
        .CO(\CARRYB[20][2] ), .S(\SUMB[20][2] ) );
  FA_X1 S2_20_3 ( .A(\ab[20][3] ), .B(\CARRYB[19][3] ), .CI(\SUMB[19][4] ), 
        .CO(\CARRYB[20][3] ), .S(\SUMB[20][3] ) );
  FA_X1 S2_20_4 ( .A(\ab[20][4] ), .B(\CARRYB[19][4] ), .CI(\SUMB[19][5] ), 
        .CO(\CARRYB[20][4] ), .S(\SUMB[20][4] ) );
  FA_X1 S2_20_5 ( .A(\ab[20][5] ), .B(\CARRYB[19][5] ), .CI(\SUMB[19][6] ), 
        .CO(\CARRYB[20][5] ), .S(\SUMB[20][5] ) );
  FA_X1 S2_20_6 ( .A(\ab[20][6] ), .B(\CARRYB[19][6] ), .CI(\SUMB[19][7] ), 
        .CO(\CARRYB[20][6] ), .S(\SUMB[20][6] ) );
  FA_X1 S2_20_7 ( .A(\ab[20][7] ), .B(\CARRYB[19][7] ), .CI(\SUMB[19][8] ), 
        .CO(\CARRYB[20][7] ), .S(\SUMB[20][7] ) );
  FA_X1 S2_20_8 ( .A(\ab[20][8] ), .B(\CARRYB[19][8] ), .CI(\SUMB[19][9] ), 
        .CO(\CARRYB[20][8] ), .S(\SUMB[20][8] ) );
  FA_X1 S2_20_9 ( .A(\ab[20][9] ), .B(\CARRYB[19][9] ), .CI(\SUMB[19][10] ), 
        .CO(\CARRYB[20][9] ), .S(\SUMB[20][9] ) );
  FA_X1 S2_20_10 ( .A(\ab[20][10] ), .B(\CARRYB[19][10] ), .CI(\SUMB[19][11] ), 
        .CO(\CARRYB[20][10] ), .S(\SUMB[20][10] ) );
  FA_X1 S2_20_11 ( .A(\ab[20][11] ), .B(\CARRYB[19][11] ), .CI(\SUMB[19][12] ), 
        .CO(\CARRYB[20][11] ), .S(\SUMB[20][11] ) );
  FA_X1 S2_20_12 ( .A(\ab[20][12] ), .B(\CARRYB[19][12] ), .CI(\SUMB[19][13] ), 
        .CO(\CARRYB[20][12] ), .S(\SUMB[20][12] ) );
  FA_X1 S2_20_13 ( .A(\ab[20][13] ), .B(\CARRYB[19][13] ), .CI(\SUMB[19][14] ), 
        .CO(\CARRYB[20][13] ), .S(\SUMB[20][13] ) );
  FA_X1 S2_20_14 ( .A(\ab[20][14] ), .B(\CARRYB[19][14] ), .CI(\SUMB[19][15] ), 
        .CO(\CARRYB[20][14] ), .S(\SUMB[20][14] ) );
  FA_X1 S2_20_15 ( .A(\CARRYB[19][15] ), .B(\ab[20][15] ), .CI(\SUMB[19][16] ), 
        .CO(\CARRYB[20][15] ), .S(\SUMB[20][15] ) );
  FA_X1 S2_20_16 ( .A(\ab[20][16] ), .B(\CARRYB[19][16] ), .CI(\SUMB[19][17] ), 
        .CO(\CARRYB[20][16] ), .S(\SUMB[20][16] ) );
  FA_X1 S2_20_17 ( .A(\ab[20][17] ), .B(\CARRYB[19][17] ), .CI(\SUMB[19][18] ), 
        .CO(\CARRYB[20][17] ), .S(\SUMB[20][17] ) );
  FA_X1 S2_20_18 ( .A(\ab[20][18] ), .B(\CARRYB[19][18] ), .CI(\SUMB[19][19] ), 
        .CO(\CARRYB[20][18] ), .S(\SUMB[20][18] ) );
  FA_X1 S2_20_19 ( .A(\ab[20][19] ), .B(\CARRYB[19][19] ), .CI(\SUMB[19][20] ), 
        .CO(\CARRYB[20][19] ), .S(\SUMB[20][19] ) );
  FA_X1 S2_20_20 ( .A(\ab[20][20] ), .B(\CARRYB[19][20] ), .CI(\SUMB[19][21] ), 
        .CO(\CARRYB[20][20] ), .S(\SUMB[20][20] ) );
  FA_X1 S2_20_21 ( .A(\ab[20][21] ), .B(\CARRYB[19][21] ), .CI(\SUMB[19][22] ), 
        .CO(\CARRYB[20][21] ), .S(\SUMB[20][21] ) );
  FA_X1 S2_20_22 ( .A(\ab[20][22] ), .B(\CARRYB[19][22] ), .CI(\SUMB[19][23] ), 
        .CO(\CARRYB[20][22] ), .S(\SUMB[20][22] ) );
  FA_X1 S2_20_23 ( .A(\ab[20][23] ), .B(\CARRYB[19][23] ), .CI(\SUMB[19][24] ), 
        .CO(\CARRYB[20][23] ), .S(\SUMB[20][23] ) );
  FA_X1 S2_20_24 ( .A(\ab[20][24] ), .B(\CARRYB[19][24] ), .CI(\SUMB[19][25] ), 
        .CO(\CARRYB[20][24] ), .S(\SUMB[20][24] ) );
  FA_X1 S2_20_25 ( .A(\ab[20][25] ), .B(\CARRYB[19][25] ), .CI(\SUMB[19][26] ), 
        .CO(\CARRYB[20][25] ), .S(\SUMB[20][25] ) );
  FA_X1 S2_20_26 ( .A(\ab[20][26] ), .B(\CARRYB[19][26] ), .CI(\SUMB[19][27] ), 
        .CO(\CARRYB[20][26] ), .S(\SUMB[20][26] ) );
  FA_X1 S2_20_27 ( .A(\ab[20][27] ), .B(\CARRYB[19][27] ), .CI(\SUMB[19][28] ), 
        .CO(\CARRYB[20][27] ), .S(\SUMB[20][27] ) );
  FA_X1 S2_20_28 ( .A(\ab[20][28] ), .B(\CARRYB[19][28] ), .CI(\SUMB[19][29] ), 
        .CO(\CARRYB[20][28] ), .S(\SUMB[20][28] ) );
  FA_X1 S2_20_29 ( .A(\ab[20][29] ), .B(\CARRYB[19][29] ), .CI(\SUMB[19][30] ), 
        .CO(\CARRYB[20][29] ), .S(\SUMB[20][29] ) );
  FA_X1 S3_20_30 ( .A(\ab[20][30] ), .B(\CARRYB[19][30] ), .CI(\ab[19][31] ), 
        .CO(\CARRYB[20][30] ), .S(\SUMB[20][30] ) );
  FA_X1 S1_19_0 ( .A(\ab[19][0] ), .B(\CARRYB[18][0] ), .CI(\SUMB[18][1] ), 
        .CO(\CARRYB[19][0] ), .S(\A1[17] ) );
  FA_X1 S2_19_1 ( .A(\ab[19][1] ), .B(\CARRYB[18][1] ), .CI(\SUMB[18][2] ), 
        .CO(\CARRYB[19][1] ), .S(\SUMB[19][1] ) );
  FA_X1 S2_19_2 ( .A(\ab[19][2] ), .B(\CARRYB[18][2] ), .CI(\SUMB[18][3] ), 
        .CO(\CARRYB[19][2] ), .S(\SUMB[19][2] ) );
  FA_X1 S2_19_3 ( .A(\ab[19][3] ), .B(\CARRYB[18][3] ), .CI(\SUMB[18][4] ), 
        .CO(\CARRYB[19][3] ), .S(\SUMB[19][3] ) );
  FA_X1 S2_19_4 ( .A(\ab[19][4] ), .B(\CARRYB[18][4] ), .CI(\SUMB[18][5] ), 
        .CO(\CARRYB[19][4] ), .S(\SUMB[19][4] ) );
  FA_X1 S2_19_5 ( .A(\ab[19][5] ), .B(\CARRYB[18][5] ), .CI(\SUMB[18][6] ), 
        .CO(\CARRYB[19][5] ), .S(\SUMB[19][5] ) );
  FA_X1 S2_19_6 ( .A(\ab[19][6] ), .B(\CARRYB[18][6] ), .CI(\SUMB[18][7] ), 
        .CO(\CARRYB[19][6] ), .S(\SUMB[19][6] ) );
  FA_X1 S2_19_7 ( .A(\ab[19][7] ), .B(\CARRYB[18][7] ), .CI(\SUMB[18][8] ), 
        .CO(\CARRYB[19][7] ), .S(\SUMB[19][7] ) );
  FA_X1 S2_19_8 ( .A(\ab[19][8] ), .B(\CARRYB[18][8] ), .CI(\SUMB[18][9] ), 
        .CO(\CARRYB[19][8] ), .S(\SUMB[19][8] ) );
  FA_X1 S2_19_9 ( .A(\ab[19][9] ), .B(\CARRYB[18][9] ), .CI(\SUMB[18][10] ), 
        .CO(\CARRYB[19][9] ), .S(\SUMB[19][9] ) );
  FA_X1 S2_19_10 ( .A(\ab[19][10] ), .B(\CARRYB[18][10] ), .CI(\SUMB[18][11] ), 
        .CO(\CARRYB[19][10] ), .S(\SUMB[19][10] ) );
  FA_X1 S2_19_11 ( .A(\ab[19][11] ), .B(\CARRYB[18][11] ), .CI(\SUMB[18][12] ), 
        .CO(\CARRYB[19][11] ), .S(\SUMB[19][11] ) );
  FA_X1 S2_19_12 ( .A(\ab[19][12] ), .B(\CARRYB[18][12] ), .CI(\SUMB[18][13] ), 
        .CO(\CARRYB[19][12] ), .S(\SUMB[19][12] ) );
  FA_X1 S2_19_13 ( .A(\ab[19][13] ), .B(\CARRYB[18][13] ), .CI(\SUMB[18][14] ), 
        .CO(\CARRYB[19][13] ), .S(\SUMB[19][13] ) );
  FA_X1 S2_19_14 ( .A(\ab[19][14] ), .B(\CARRYB[18][14] ), .CI(\SUMB[18][15] ), 
        .CO(\CARRYB[19][14] ), .S(\SUMB[19][14] ) );
  FA_X1 S2_19_15 ( .A(\ab[19][15] ), .B(\CARRYB[18][15] ), .CI(\SUMB[18][16] ), 
        .CO(\CARRYB[19][15] ), .S(\SUMB[19][15] ) );
  FA_X1 S2_19_16 ( .A(\ab[19][16] ), .B(\CARRYB[18][16] ), .CI(\SUMB[18][17] ), 
        .CO(\CARRYB[19][16] ), .S(\SUMB[19][16] ) );
  FA_X1 S2_19_17 ( .A(\ab[19][17] ), .B(\CARRYB[18][17] ), .CI(\SUMB[18][18] ), 
        .CO(\CARRYB[19][17] ), .S(\SUMB[19][17] ) );
  FA_X1 S2_19_18 ( .A(\ab[19][18] ), .B(\CARRYB[18][18] ), .CI(\SUMB[18][19] ), 
        .CO(\CARRYB[19][18] ), .S(\SUMB[19][18] ) );
  FA_X1 S2_19_19 ( .A(\ab[19][19] ), .B(\CARRYB[18][19] ), .CI(\SUMB[18][20] ), 
        .CO(\CARRYB[19][19] ), .S(\SUMB[19][19] ) );
  FA_X1 S2_19_20 ( .A(\ab[19][20] ), .B(\CARRYB[18][20] ), .CI(\SUMB[18][21] ), 
        .CO(\CARRYB[19][20] ), .S(\SUMB[19][20] ) );
  FA_X1 S2_19_21 ( .A(\ab[19][21] ), .B(\CARRYB[18][21] ), .CI(\SUMB[18][22] ), 
        .CO(\CARRYB[19][21] ), .S(\SUMB[19][21] ) );
  FA_X1 S2_19_22 ( .A(\ab[19][22] ), .B(\CARRYB[18][22] ), .CI(\SUMB[18][23] ), 
        .CO(\CARRYB[19][22] ), .S(\SUMB[19][22] ) );
  FA_X1 S2_19_23 ( .A(\ab[19][23] ), .B(\CARRYB[18][23] ), .CI(\SUMB[18][24] ), 
        .CO(\CARRYB[19][23] ), .S(\SUMB[19][23] ) );
  FA_X1 S2_19_24 ( .A(\ab[19][24] ), .B(\CARRYB[18][24] ), .CI(\SUMB[18][25] ), 
        .CO(\CARRYB[19][24] ), .S(\SUMB[19][24] ) );
  FA_X1 S2_19_25 ( .A(\ab[19][25] ), .B(\CARRYB[18][25] ), .CI(\SUMB[18][26] ), 
        .CO(\CARRYB[19][25] ), .S(\SUMB[19][25] ) );
  FA_X1 S2_19_26 ( .A(\ab[19][26] ), .B(\CARRYB[18][26] ), .CI(\SUMB[18][27] ), 
        .CO(\CARRYB[19][26] ), .S(\SUMB[19][26] ) );
  FA_X1 S2_19_27 ( .A(\ab[19][27] ), .B(\CARRYB[18][27] ), .CI(\SUMB[18][28] ), 
        .CO(\CARRYB[19][27] ), .S(\SUMB[19][27] ) );
  FA_X1 S2_19_28 ( .A(\ab[19][28] ), .B(\CARRYB[18][28] ), .CI(\SUMB[18][29] ), 
        .CO(\CARRYB[19][28] ), .S(\SUMB[19][28] ) );
  FA_X1 S2_19_29 ( .A(\ab[19][29] ), .B(\CARRYB[18][29] ), .CI(\SUMB[18][30] ), 
        .CO(\CARRYB[19][29] ), .S(\SUMB[19][29] ) );
  FA_X1 S3_19_30 ( .A(\ab[19][30] ), .B(\CARRYB[18][30] ), .CI(\ab[18][31] ), 
        .CO(\CARRYB[19][30] ), .S(\SUMB[19][30] ) );
  FA_X1 S1_18_0 ( .A(\ab[18][0] ), .B(\CARRYB[17][0] ), .CI(\SUMB[17][1] ), 
        .CO(\CARRYB[18][0] ), .S(\A1[16] ) );
  FA_X1 S2_18_1 ( .A(\ab[18][1] ), .B(\CARRYB[17][1] ), .CI(\SUMB[17][2] ), 
        .CO(\CARRYB[18][1] ), .S(\SUMB[18][1] ) );
  FA_X1 S2_18_2 ( .A(\ab[18][2] ), .B(\CARRYB[17][2] ), .CI(\SUMB[17][3] ), 
        .CO(\CARRYB[18][2] ), .S(\SUMB[18][2] ) );
  FA_X1 S2_18_3 ( .A(\ab[18][3] ), .B(\CARRYB[17][3] ), .CI(\SUMB[17][4] ), 
        .CO(\CARRYB[18][3] ), .S(\SUMB[18][3] ) );
  FA_X1 S2_18_4 ( .A(\ab[18][4] ), .B(\CARRYB[17][4] ), .CI(\SUMB[17][5] ), 
        .CO(\CARRYB[18][4] ), .S(\SUMB[18][4] ) );
  FA_X1 S2_18_5 ( .A(\ab[18][5] ), .B(\CARRYB[17][5] ), .CI(\SUMB[17][6] ), 
        .CO(\CARRYB[18][5] ), .S(\SUMB[18][5] ) );
  FA_X1 S2_18_6 ( .A(\ab[18][6] ), .B(\CARRYB[17][6] ), .CI(\SUMB[17][7] ), 
        .CO(\CARRYB[18][6] ), .S(\SUMB[18][6] ) );
  FA_X1 S2_18_7 ( .A(\ab[18][7] ), .B(\CARRYB[17][7] ), .CI(\SUMB[17][8] ), 
        .CO(\CARRYB[18][7] ), .S(\SUMB[18][7] ) );
  FA_X1 S2_18_8 ( .A(\ab[18][8] ), .B(\CARRYB[17][8] ), .CI(\SUMB[17][9] ), 
        .CO(\CARRYB[18][8] ), .S(\SUMB[18][8] ) );
  FA_X1 S2_18_9 ( .A(\ab[18][9] ), .B(\CARRYB[17][9] ), .CI(\SUMB[17][10] ), 
        .CO(\CARRYB[18][9] ), .S(\SUMB[18][9] ) );
  FA_X1 S2_18_10 ( .A(\ab[18][10] ), .B(\CARRYB[17][10] ), .CI(\SUMB[17][11] ), 
        .CO(\CARRYB[18][10] ), .S(\SUMB[18][10] ) );
  FA_X1 S2_18_11 ( .A(\ab[18][11] ), .B(\CARRYB[17][11] ), .CI(\SUMB[17][12] ), 
        .CO(\CARRYB[18][11] ), .S(\SUMB[18][11] ) );
  FA_X1 S2_18_12 ( .A(\ab[18][12] ), .B(\CARRYB[17][12] ), .CI(\SUMB[17][13] ), 
        .CO(\CARRYB[18][12] ), .S(\SUMB[18][12] ) );
  FA_X1 S2_18_13 ( .A(\ab[18][13] ), .B(\CARRYB[17][13] ), .CI(\SUMB[17][14] ), 
        .CO(\CARRYB[18][13] ), .S(\SUMB[18][13] ) );
  FA_X1 S2_18_14 ( .A(\ab[18][14] ), .B(\CARRYB[17][14] ), .CI(\SUMB[17][15] ), 
        .CO(\CARRYB[18][14] ), .S(\SUMB[18][14] ) );
  FA_X1 S2_18_15 ( .A(\ab[18][15] ), .B(\CARRYB[17][15] ), .CI(\SUMB[17][16] ), 
        .CO(\CARRYB[18][15] ), .S(\SUMB[18][15] ) );
  FA_X1 S2_18_16 ( .A(\ab[18][16] ), .B(\CARRYB[17][16] ), .CI(\SUMB[17][17] ), 
        .CO(\CARRYB[18][16] ), .S(\SUMB[18][16] ) );
  FA_X1 S2_18_17 ( .A(\ab[18][17] ), .B(\CARRYB[17][17] ), .CI(\SUMB[17][18] ), 
        .CO(\CARRYB[18][17] ), .S(\SUMB[18][17] ) );
  FA_X1 S2_18_18 ( .A(\ab[18][18] ), .B(\CARRYB[17][18] ), .CI(\SUMB[17][19] ), 
        .CO(\CARRYB[18][18] ), .S(\SUMB[18][18] ) );
  FA_X1 S2_18_19 ( .A(\ab[18][19] ), .B(\CARRYB[17][19] ), .CI(\SUMB[17][20] ), 
        .CO(\CARRYB[18][19] ), .S(\SUMB[18][19] ) );
  FA_X1 S2_18_20 ( .A(\ab[18][20] ), .B(\CARRYB[17][20] ), .CI(\SUMB[17][21] ), 
        .CO(\CARRYB[18][20] ), .S(\SUMB[18][20] ) );
  FA_X1 S2_18_21 ( .A(\ab[18][21] ), .B(\CARRYB[17][21] ), .CI(\SUMB[17][22] ), 
        .CO(\CARRYB[18][21] ), .S(\SUMB[18][21] ) );
  FA_X1 S2_18_22 ( .A(\ab[18][22] ), .B(\CARRYB[17][22] ), .CI(\SUMB[17][23] ), 
        .CO(\CARRYB[18][22] ), .S(\SUMB[18][22] ) );
  FA_X1 S2_18_23 ( .A(\ab[18][23] ), .B(\CARRYB[17][23] ), .CI(\SUMB[17][24] ), 
        .CO(\CARRYB[18][23] ), .S(\SUMB[18][23] ) );
  FA_X1 S2_18_24 ( .A(\ab[18][24] ), .B(\CARRYB[17][24] ), .CI(\SUMB[17][25] ), 
        .CO(\CARRYB[18][24] ), .S(\SUMB[18][24] ) );
  FA_X1 S2_18_25 ( .A(\ab[18][25] ), .B(\CARRYB[17][25] ), .CI(\SUMB[17][26] ), 
        .CO(\CARRYB[18][25] ), .S(\SUMB[18][25] ) );
  FA_X1 S2_18_26 ( .A(\ab[18][26] ), .B(\CARRYB[17][26] ), .CI(\SUMB[17][27] ), 
        .CO(\CARRYB[18][26] ), .S(\SUMB[18][26] ) );
  FA_X1 S2_18_27 ( .A(\ab[18][27] ), .B(\CARRYB[17][27] ), .CI(\SUMB[17][28] ), 
        .CO(\CARRYB[18][27] ), .S(\SUMB[18][27] ) );
  FA_X1 S2_18_28 ( .A(\ab[18][28] ), .B(\CARRYB[17][28] ), .CI(\SUMB[17][29] ), 
        .CO(\CARRYB[18][28] ), .S(\SUMB[18][28] ) );
  FA_X1 S2_18_29 ( .A(\ab[18][29] ), .B(\CARRYB[17][29] ), .CI(\SUMB[17][30] ), 
        .CO(\CARRYB[18][29] ), .S(\SUMB[18][29] ) );
  FA_X1 S3_18_30 ( .A(\ab[18][30] ), .B(\CARRYB[17][30] ), .CI(\ab[17][31] ), 
        .CO(\CARRYB[18][30] ), .S(\SUMB[18][30] ) );
  FA_X1 S1_17_0 ( .A(\ab[17][0] ), .B(\CARRYB[16][0] ), .CI(\SUMB[16][1] ), 
        .CO(\CARRYB[17][0] ), .S(\A1[15] ) );
  FA_X1 S2_17_1 ( .A(\ab[17][1] ), .B(\CARRYB[16][1] ), .CI(\SUMB[16][2] ), 
        .CO(\CARRYB[17][1] ), .S(\SUMB[17][1] ) );
  FA_X1 S2_17_2 ( .A(\ab[17][2] ), .B(\CARRYB[16][2] ), .CI(\SUMB[16][3] ), 
        .CO(\CARRYB[17][2] ), .S(\SUMB[17][2] ) );
  FA_X1 S2_17_3 ( .A(\ab[17][3] ), .B(\CARRYB[16][3] ), .CI(\SUMB[16][4] ), 
        .CO(\CARRYB[17][3] ), .S(\SUMB[17][3] ) );
  FA_X1 S2_17_4 ( .A(\ab[17][4] ), .B(\CARRYB[16][4] ), .CI(\SUMB[16][5] ), 
        .CO(\CARRYB[17][4] ), .S(\SUMB[17][4] ) );
  FA_X1 S2_17_5 ( .A(\ab[17][5] ), .B(\CARRYB[16][5] ), .CI(\SUMB[16][6] ), 
        .CO(\CARRYB[17][5] ), .S(\SUMB[17][5] ) );
  FA_X1 S2_17_6 ( .A(\ab[17][6] ), .B(\CARRYB[16][6] ), .CI(\SUMB[16][7] ), 
        .CO(\CARRYB[17][6] ), .S(\SUMB[17][6] ) );
  FA_X1 S2_17_7 ( .A(\ab[17][7] ), .B(\CARRYB[16][7] ), .CI(\SUMB[16][8] ), 
        .CO(\CARRYB[17][7] ), .S(\SUMB[17][7] ) );
  FA_X1 S2_17_8 ( .A(\ab[17][8] ), .B(\CARRYB[16][8] ), .CI(\SUMB[16][9] ), 
        .CO(\CARRYB[17][8] ), .S(\SUMB[17][8] ) );
  FA_X1 S2_17_9 ( .A(\ab[17][9] ), .B(\CARRYB[16][9] ), .CI(\SUMB[16][10] ), 
        .CO(\CARRYB[17][9] ), .S(\SUMB[17][9] ) );
  FA_X1 S2_17_10 ( .A(\ab[17][10] ), .B(\CARRYB[16][10] ), .CI(\SUMB[16][11] ), 
        .CO(\CARRYB[17][10] ), .S(\SUMB[17][10] ) );
  FA_X1 S2_17_11 ( .A(\ab[17][11] ), .B(\CARRYB[16][11] ), .CI(\SUMB[16][12] ), 
        .CO(\CARRYB[17][11] ), .S(\SUMB[17][11] ) );
  FA_X1 S2_17_12 ( .A(\ab[17][12] ), .B(\CARRYB[16][12] ), .CI(\SUMB[16][13] ), 
        .CO(\CARRYB[17][12] ), .S(\SUMB[17][12] ) );
  FA_X1 S2_17_13 ( .A(\ab[17][13] ), .B(\CARRYB[16][13] ), .CI(\SUMB[16][14] ), 
        .CO(\CARRYB[17][13] ), .S(\SUMB[17][13] ) );
  FA_X1 S2_17_14 ( .A(\ab[17][14] ), .B(\CARRYB[16][14] ), .CI(\SUMB[16][15] ), 
        .CO(\CARRYB[17][14] ), .S(\SUMB[17][14] ) );
  FA_X1 S2_17_15 ( .A(\ab[17][15] ), .B(\CARRYB[16][15] ), .CI(\SUMB[16][16] ), 
        .CO(\CARRYB[17][15] ), .S(\SUMB[17][15] ) );
  FA_X1 S2_17_16 ( .A(\ab[17][16] ), .B(\CARRYB[16][16] ), .CI(\SUMB[16][17] ), 
        .CO(\CARRYB[17][16] ), .S(\SUMB[17][16] ) );
  FA_X1 S2_17_17 ( .A(\CARRYB[16][17] ), .B(\ab[17][17] ), .CI(\SUMB[16][18] ), 
        .CO(\CARRYB[17][17] ), .S(\SUMB[17][17] ) );
  FA_X1 S2_17_18 ( .A(\ab[17][18] ), .B(\CARRYB[16][18] ), .CI(\SUMB[16][19] ), 
        .CO(\CARRYB[17][18] ), .S(\SUMB[17][18] ) );
  FA_X1 S2_17_19 ( .A(\ab[17][19] ), .B(\CARRYB[16][19] ), .CI(\SUMB[16][20] ), 
        .CO(\CARRYB[17][19] ), .S(\SUMB[17][19] ) );
  FA_X1 S2_17_20 ( .A(\ab[17][20] ), .B(\CARRYB[16][20] ), .CI(\SUMB[16][21] ), 
        .CO(\CARRYB[17][20] ), .S(\SUMB[17][20] ) );
  FA_X1 S2_17_21 ( .A(\ab[17][21] ), .B(\CARRYB[16][21] ), .CI(\SUMB[16][22] ), 
        .CO(\CARRYB[17][21] ), .S(\SUMB[17][21] ) );
  FA_X1 S2_17_22 ( .A(\ab[17][22] ), .B(\CARRYB[16][22] ), .CI(\SUMB[16][23] ), 
        .CO(\CARRYB[17][22] ), .S(\SUMB[17][22] ) );
  FA_X1 S2_17_23 ( .A(\ab[17][23] ), .B(\CARRYB[16][23] ), .CI(\SUMB[16][24] ), 
        .CO(\CARRYB[17][23] ), .S(\SUMB[17][23] ) );
  FA_X1 S2_17_24 ( .A(\ab[17][24] ), .B(\CARRYB[16][24] ), .CI(\SUMB[16][25] ), 
        .CO(\CARRYB[17][24] ), .S(\SUMB[17][24] ) );
  FA_X1 S2_17_25 ( .A(\ab[17][25] ), .B(\CARRYB[16][25] ), .CI(\SUMB[16][26] ), 
        .CO(\CARRYB[17][25] ), .S(\SUMB[17][25] ) );
  FA_X1 S2_17_26 ( .A(\ab[17][26] ), .B(\CARRYB[16][26] ), .CI(\SUMB[16][27] ), 
        .CO(\CARRYB[17][26] ), .S(\SUMB[17][26] ) );
  FA_X1 S2_17_27 ( .A(\ab[17][27] ), .B(\CARRYB[16][27] ), .CI(\SUMB[16][28] ), 
        .CO(\CARRYB[17][27] ), .S(\SUMB[17][27] ) );
  FA_X1 S2_17_28 ( .A(\ab[17][28] ), .B(\CARRYB[16][28] ), .CI(\SUMB[16][29] ), 
        .CO(\CARRYB[17][28] ), .S(\SUMB[17][28] ) );
  FA_X1 S2_17_29 ( .A(\ab[17][29] ), .B(\CARRYB[16][29] ), .CI(\SUMB[16][30] ), 
        .CO(\CARRYB[17][29] ), .S(\SUMB[17][29] ) );
  FA_X1 S3_17_30 ( .A(\ab[17][30] ), .B(\CARRYB[16][30] ), .CI(\ab[16][31] ), 
        .CO(\CARRYB[17][30] ), .S(\SUMB[17][30] ) );
  FA_X1 S1_16_0 ( .A(\ab[16][0] ), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), 
        .CO(\CARRYB[16][0] ), .S(\A1[14] ) );
  FA_X1 S2_16_1 ( .A(\ab[16][1] ), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), 
        .CO(\CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FA_X1 S2_16_2 ( .A(\ab[16][2] ), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), 
        .CO(\CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FA_X1 S2_16_3 ( .A(\ab[16][3] ), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), 
        .CO(\CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FA_X1 S2_16_4 ( .A(\ab[16][4] ), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), 
        .CO(\CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FA_X1 S2_16_5 ( .A(\ab[16][5] ), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), 
        .CO(\CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FA_X1 S2_16_6 ( .A(\ab[16][6] ), .B(\CARRYB[15][6] ), .CI(\SUMB[15][7] ), 
        .CO(\CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FA_X1 S2_16_7 ( .A(\ab[16][7] ), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), 
        .CO(\CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FA_X1 S2_16_8 ( .A(\ab[16][8] ), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), 
        .CO(\CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FA_X1 S2_16_9 ( .A(\ab[16][9] ), .B(\CARRYB[15][9] ), .CI(\SUMB[15][10] ), 
        .CO(\CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FA_X1 S2_16_10 ( .A(\ab[16][10] ), .B(\CARRYB[15][10] ), .CI(\SUMB[15][11] ), 
        .CO(\CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FA_X1 S2_16_11 ( .A(\ab[16][11] ), .B(\CARRYB[15][11] ), .CI(\SUMB[15][12] ), 
        .CO(\CARRYB[16][11] ), .S(\SUMB[16][11] ) );
  FA_X1 S2_16_12 ( .A(\ab[16][12] ), .B(\CARRYB[15][12] ), .CI(\SUMB[15][13] ), 
        .CO(\CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FA_X1 S2_16_13 ( .A(\ab[16][13] ), .B(\CARRYB[15][13] ), .CI(\SUMB[15][14] ), 
        .CO(\CARRYB[16][13] ), .S(\SUMB[16][13] ) );
  FA_X1 S2_16_14 ( .A(\ab[16][14] ), .B(\CARRYB[15][14] ), .CI(\SUMB[15][15] ), 
        .CO(\CARRYB[16][14] ), .S(\SUMB[16][14] ) );
  FA_X1 S2_16_15 ( .A(\ab[16][15] ), .B(\CARRYB[15][15] ), .CI(\SUMB[15][16] ), 
        .CO(\CARRYB[16][15] ), .S(\SUMB[16][15] ) );
  FA_X1 S2_16_16 ( .A(\ab[16][16] ), .B(\CARRYB[15][16] ), .CI(\SUMB[15][17] ), 
        .CO(\CARRYB[16][16] ), .S(\SUMB[16][16] ) );
  FA_X1 S2_16_17 ( .A(\ab[16][17] ), .B(\CARRYB[15][17] ), .CI(\SUMB[15][18] ), 
        .CO(\CARRYB[16][17] ), .S(\SUMB[16][17] ) );
  FA_X1 S2_16_18 ( .A(\ab[16][18] ), .B(\CARRYB[15][18] ), .CI(\SUMB[15][19] ), 
        .CO(\CARRYB[16][18] ), .S(\SUMB[16][18] ) );
  FA_X1 S2_16_19 ( .A(\ab[16][19] ), .B(\CARRYB[15][19] ), .CI(\SUMB[15][20] ), 
        .CO(\CARRYB[16][19] ), .S(\SUMB[16][19] ) );
  FA_X1 S2_16_20 ( .A(\ab[16][20] ), .B(\CARRYB[15][20] ), .CI(\SUMB[15][21] ), 
        .CO(\CARRYB[16][20] ), .S(\SUMB[16][20] ) );
  FA_X1 S2_16_21 ( .A(\ab[16][21] ), .B(\CARRYB[15][21] ), .CI(\SUMB[15][22] ), 
        .CO(\CARRYB[16][21] ), .S(\SUMB[16][21] ) );
  FA_X1 S2_16_22 ( .A(\ab[16][22] ), .B(\CARRYB[15][22] ), .CI(\SUMB[15][23] ), 
        .CO(\CARRYB[16][22] ), .S(\SUMB[16][22] ) );
  FA_X1 S2_16_23 ( .A(\ab[16][23] ), .B(\CARRYB[15][23] ), .CI(\SUMB[15][24] ), 
        .CO(\CARRYB[16][23] ), .S(\SUMB[16][23] ) );
  FA_X1 S2_16_24 ( .A(\ab[16][24] ), .B(\CARRYB[15][24] ), .CI(\SUMB[15][25] ), 
        .CO(\CARRYB[16][24] ), .S(\SUMB[16][24] ) );
  FA_X1 S2_16_25 ( .A(\ab[16][25] ), .B(\CARRYB[15][25] ), .CI(\SUMB[15][26] ), 
        .CO(\CARRYB[16][25] ), .S(\SUMB[16][25] ) );
  FA_X1 S2_16_26 ( .A(\ab[16][26] ), .B(\CARRYB[15][26] ), .CI(\SUMB[15][27] ), 
        .CO(\CARRYB[16][26] ), .S(\SUMB[16][26] ) );
  FA_X1 S2_16_27 ( .A(\ab[16][27] ), .B(\CARRYB[15][27] ), .CI(\SUMB[15][28] ), 
        .CO(\CARRYB[16][27] ), .S(\SUMB[16][27] ) );
  FA_X1 S2_16_28 ( .A(\ab[16][28] ), .B(\CARRYB[15][28] ), .CI(\SUMB[15][29] ), 
        .CO(\CARRYB[16][28] ), .S(\SUMB[16][28] ) );
  FA_X1 S2_16_29 ( .A(\ab[16][29] ), .B(\CARRYB[15][29] ), .CI(\SUMB[15][30] ), 
        .CO(\CARRYB[16][29] ), .S(\SUMB[16][29] ) );
  FA_X1 S3_16_30 ( .A(\ab[16][30] ), .B(\CARRYB[15][30] ), .CI(\ab[15][31] ), 
        .CO(\CARRYB[16][30] ), .S(\SUMB[16][30] ) );
  FA_X1 S1_15_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), 
        .CO(\CARRYB[15][0] ), .S(\A1[13] ) );
  FA_X1 S2_15_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), 
        .CO(\CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA_X1 S2_15_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), 
        .CO(\CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA_X1 S2_15_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), 
        .CO(\CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA_X1 S2_15_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), 
        .CO(\CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA_X1 S2_15_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), 
        .CO(\CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA_X1 S2_15_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), 
        .CO(\CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA_X1 S2_15_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), 
        .CO(\CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA_X1 S2_15_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), 
        .CO(\CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA_X1 S2_15_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), 
        .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA_X1 S2_15_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA_X1 S2_15_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA_X1 S2_15_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA_X1 S2_15_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA_X1 S2_15_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\SUMB[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA_X1 S2_15_15 ( .A(\ab[15][15] ), .B(\CARRYB[14][15] ), .CI(\SUMB[14][16] ), 
        .CO(\CARRYB[15][15] ), .S(\SUMB[15][15] ) );
  FA_X1 S2_15_16 ( .A(\CARRYB[14][16] ), .B(\ab[15][16] ), .CI(\SUMB[14][17] ), 
        .CO(\CARRYB[15][16] ), .S(\SUMB[15][16] ) );
  FA_X1 S2_15_17 ( .A(\CARRYB[14][17] ), .B(\ab[15][17] ), .CI(\SUMB[14][18] ), 
        .CO(\CARRYB[15][17] ), .S(\SUMB[15][17] ) );
  FA_X1 S2_15_18 ( .A(\ab[15][18] ), .B(\CARRYB[14][18] ), .CI(\SUMB[14][19] ), 
        .CO(\CARRYB[15][18] ), .S(\SUMB[15][18] ) );
  FA_X1 S2_15_19 ( .A(\CARRYB[14][19] ), .B(\ab[15][19] ), .CI(\SUMB[14][20] ), 
        .CO(\CARRYB[15][19] ), .S(\SUMB[15][19] ) );
  FA_X1 S2_15_20 ( .A(\ab[15][20] ), .B(\CARRYB[14][20] ), .CI(\SUMB[14][21] ), 
        .CO(\CARRYB[15][20] ), .S(\SUMB[15][20] ) );
  FA_X1 S2_15_21 ( .A(\ab[15][21] ), .B(\CARRYB[14][21] ), .CI(\SUMB[14][22] ), 
        .CO(\CARRYB[15][21] ), .S(\SUMB[15][21] ) );
  FA_X1 S2_15_22 ( .A(\ab[15][22] ), .B(\CARRYB[14][22] ), .CI(\SUMB[14][23] ), 
        .CO(\CARRYB[15][22] ), .S(\SUMB[15][22] ) );
  FA_X1 S2_15_23 ( .A(\ab[15][23] ), .B(\CARRYB[14][23] ), .CI(\SUMB[14][24] ), 
        .CO(\CARRYB[15][23] ), .S(\SUMB[15][23] ) );
  FA_X1 S2_15_24 ( .A(\ab[15][24] ), .B(\CARRYB[14][24] ), .CI(\SUMB[14][25] ), 
        .CO(\CARRYB[15][24] ), .S(\SUMB[15][24] ) );
  FA_X1 S2_15_25 ( .A(\ab[15][25] ), .B(\CARRYB[14][25] ), .CI(\SUMB[14][26] ), 
        .CO(\CARRYB[15][25] ), .S(\SUMB[15][25] ) );
  FA_X1 S2_15_26 ( .A(\ab[15][26] ), .B(\CARRYB[14][26] ), .CI(\SUMB[14][27] ), 
        .CO(\CARRYB[15][26] ), .S(\SUMB[15][26] ) );
  FA_X1 S2_15_27 ( .A(\ab[15][27] ), .B(\CARRYB[14][27] ), .CI(\SUMB[14][28] ), 
        .CO(\CARRYB[15][27] ), .S(\SUMB[15][27] ) );
  FA_X1 S2_15_28 ( .A(\ab[15][28] ), .B(\CARRYB[14][28] ), .CI(\SUMB[14][29] ), 
        .CO(\CARRYB[15][28] ), .S(\SUMB[15][28] ) );
  FA_X1 S2_15_29 ( .A(\ab[15][29] ), .B(\CARRYB[14][29] ), .CI(\SUMB[14][30] ), 
        .CO(\CARRYB[15][29] ), .S(\SUMB[15][29] ) );
  FA_X1 S3_15_30 ( .A(\ab[15][30] ), .B(\CARRYB[14][30] ), .CI(\ab[14][31] ), 
        .CO(\CARRYB[15][30] ), .S(\SUMB[15][30] ) );
  FA_X1 S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FA_X1 S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA_X1 S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA_X1 S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA_X1 S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA_X1 S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA_X1 S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA_X1 S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA_X1 S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA_X1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA_X1 S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA_X1 S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA_X1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA_X1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA_X1 S2_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA_X1 S2_14_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(\SUMB[13][16] ), 
        .CO(\CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FA_X1 S2_14_16 ( .A(\ab[14][16] ), .B(\CARRYB[13][16] ), .CI(\SUMB[13][17] ), 
        .CO(\CARRYB[14][16] ), .S(\SUMB[14][16] ) );
  FA_X1 S2_14_17 ( .A(\ab[14][17] ), .B(\CARRYB[13][17] ), .CI(\SUMB[13][18] ), 
        .CO(\CARRYB[14][17] ), .S(\SUMB[14][17] ) );
  FA_X1 S2_14_18 ( .A(\ab[14][18] ), .B(\CARRYB[13][18] ), .CI(\SUMB[13][19] ), 
        .CO(\CARRYB[14][18] ), .S(\SUMB[14][18] ) );
  FA_X1 S2_14_19 ( .A(\CARRYB[13][19] ), .B(\ab[14][19] ), .CI(\SUMB[13][20] ), 
        .CO(\CARRYB[14][19] ), .S(\SUMB[14][19] ) );
  FA_X1 S2_14_20 ( .A(\ab[14][20] ), .B(\CARRYB[13][20] ), .CI(\SUMB[13][21] ), 
        .CO(\CARRYB[14][20] ), .S(\SUMB[14][20] ) );
  FA_X1 S2_14_21 ( .A(\ab[14][21] ), .B(\CARRYB[13][21] ), .CI(\SUMB[13][22] ), 
        .CO(\CARRYB[14][21] ), .S(\SUMB[14][21] ) );
  FA_X1 S2_14_22 ( .A(\ab[14][22] ), .B(\CARRYB[13][22] ), .CI(\SUMB[13][23] ), 
        .CO(\CARRYB[14][22] ), .S(\SUMB[14][22] ) );
  FA_X1 S2_14_23 ( .A(\ab[14][23] ), .B(\CARRYB[13][23] ), .CI(\SUMB[13][24] ), 
        .CO(\CARRYB[14][23] ), .S(\SUMB[14][23] ) );
  FA_X1 S2_14_24 ( .A(\ab[14][24] ), .B(\CARRYB[13][24] ), .CI(\SUMB[13][25] ), 
        .CO(\CARRYB[14][24] ), .S(\SUMB[14][24] ) );
  FA_X1 S2_14_25 ( .A(\ab[14][25] ), .B(\CARRYB[13][25] ), .CI(\SUMB[13][26] ), 
        .CO(\CARRYB[14][25] ), .S(\SUMB[14][25] ) );
  FA_X1 S2_14_26 ( .A(\ab[14][26] ), .B(\CARRYB[13][26] ), .CI(\SUMB[13][27] ), 
        .CO(\CARRYB[14][26] ), .S(\SUMB[14][26] ) );
  FA_X1 S2_14_27 ( .A(\ab[14][27] ), .B(\CARRYB[13][27] ), .CI(\SUMB[13][28] ), 
        .CO(\CARRYB[14][27] ), .S(\SUMB[14][27] ) );
  FA_X1 S2_14_28 ( .A(\ab[14][28] ), .B(\CARRYB[13][28] ), .CI(\SUMB[13][29] ), 
        .CO(\CARRYB[14][28] ), .S(\SUMB[14][28] ) );
  FA_X1 S2_14_29 ( .A(\ab[14][29] ), .B(\CARRYB[13][29] ), .CI(\SUMB[13][30] ), 
        .CO(\CARRYB[14][29] ), .S(\SUMB[14][29] ) );
  FA_X1 S3_14_30 ( .A(\ab[14][30] ), .B(\CARRYB[13][30] ), .CI(\ab[13][31] ), 
        .CO(\CARRYB[14][30] ), .S(\SUMB[14][30] ) );
  FA_X1 S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA_X1 S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA_X1 S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA_X1 S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA_X1 S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA_X1 S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA_X1 S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA_X1 S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA_X1 S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA_X1 S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA_X1 S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA_X1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA_X1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA_X1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA_X1 S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA_X1 S2_13_15 ( .A(\ab[13][15] ), .B(\CARRYB[12][15] ), .CI(\SUMB[12][16] ), 
        .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA_X1 S2_13_16 ( .A(\ab[13][16] ), .B(\CARRYB[12][16] ), .CI(\SUMB[12][17] ), 
        .CO(\CARRYB[13][16] ), .S(\SUMB[13][16] ) );
  FA_X1 S2_13_17 ( .A(\ab[13][17] ), .B(\CARRYB[12][17] ), .CI(\SUMB[12][18] ), 
        .CO(\CARRYB[13][17] ), .S(\SUMB[13][17] ) );
  FA_X1 S2_13_18 ( .A(\ab[13][18] ), .B(\CARRYB[12][18] ), .CI(\SUMB[12][19] ), 
        .CO(\CARRYB[13][18] ), .S(\SUMB[13][18] ) );
  FA_X1 S2_13_19 ( .A(\ab[13][19] ), .B(\CARRYB[12][19] ), .CI(\SUMB[12][20] ), 
        .CO(\CARRYB[13][19] ), .S(\SUMB[13][19] ) );
  FA_X1 S2_13_20 ( .A(\ab[13][20] ), .B(\CARRYB[12][20] ), .CI(\SUMB[12][21] ), 
        .CO(\CARRYB[13][20] ), .S(\SUMB[13][20] ) );
  FA_X1 S2_13_21 ( .A(\CARRYB[12][21] ), .B(\ab[13][21] ), .CI(\SUMB[12][22] ), 
        .CO(\CARRYB[13][21] ), .S(\SUMB[13][21] ) );
  FA_X1 S2_13_22 ( .A(\ab[13][22] ), .B(\CARRYB[12][22] ), .CI(\SUMB[12][23] ), 
        .CO(\CARRYB[13][22] ), .S(\SUMB[13][22] ) );
  FA_X1 S2_13_23 ( .A(\ab[13][23] ), .B(\CARRYB[12][23] ), .CI(\SUMB[12][24] ), 
        .CO(\CARRYB[13][23] ), .S(\SUMB[13][23] ) );
  FA_X1 S2_13_24 ( .A(\ab[13][24] ), .B(\CARRYB[12][24] ), .CI(\SUMB[12][25] ), 
        .CO(\CARRYB[13][24] ), .S(\SUMB[13][24] ) );
  FA_X1 S2_13_25 ( .A(\ab[13][25] ), .B(\CARRYB[12][25] ), .CI(\SUMB[12][26] ), 
        .CO(\CARRYB[13][25] ), .S(\SUMB[13][25] ) );
  FA_X1 S2_13_26 ( .A(\ab[13][26] ), .B(\CARRYB[12][26] ), .CI(\SUMB[12][27] ), 
        .CO(\CARRYB[13][26] ), .S(\SUMB[13][26] ) );
  FA_X1 S2_13_27 ( .A(\ab[13][27] ), .B(\CARRYB[12][27] ), .CI(\SUMB[12][28] ), 
        .CO(\CARRYB[13][27] ), .S(\SUMB[13][27] ) );
  FA_X1 S2_13_28 ( .A(\ab[13][28] ), .B(\CARRYB[12][28] ), .CI(\SUMB[12][29] ), 
        .CO(\CARRYB[13][28] ), .S(\SUMB[13][28] ) );
  FA_X1 S2_13_29 ( .A(\ab[13][29] ), .B(\CARRYB[12][29] ), .CI(\SUMB[12][30] ), 
        .CO(\CARRYB[13][29] ), .S(\SUMB[13][29] ) );
  FA_X1 S3_13_30 ( .A(\ab[13][30] ), .B(\CARRYB[12][30] ), .CI(\ab[12][31] ), 
        .CO(\CARRYB[13][30] ), .S(\SUMB[13][30] ) );
  FA_X1 S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA_X1 S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA_X1 S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA_X1 S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA_X1 S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA_X1 S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA_X1 S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA_X1 S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA_X1 S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA_X1 S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA_X1 S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA_X1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA_X1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA_X1 S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA_X1 S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA_X1 S2_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(\SUMB[11][16] ), 
        .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA_X1 S2_12_16 ( .A(\ab[12][16] ), .B(\CARRYB[11][16] ), .CI(\SUMB[11][17] ), 
        .CO(\CARRYB[12][16] ), .S(\SUMB[12][16] ) );
  FA_X1 S2_12_17 ( .A(\ab[12][17] ), .B(\CARRYB[11][17] ), .CI(\SUMB[11][18] ), 
        .CO(\CARRYB[12][17] ), .S(\SUMB[12][17] ) );
  FA_X1 S2_12_18 ( .A(\ab[12][18] ), .B(\CARRYB[11][18] ), .CI(\SUMB[11][19] ), 
        .CO(\CARRYB[12][18] ), .S(\SUMB[12][18] ) );
  FA_X1 S2_12_19 ( .A(\ab[12][19] ), .B(\CARRYB[11][19] ), .CI(\SUMB[11][20] ), 
        .CO(\CARRYB[12][19] ), .S(\SUMB[12][19] ) );
  FA_X1 S2_12_20 ( .A(\ab[12][20] ), .B(\CARRYB[11][20] ), .CI(\SUMB[11][21] ), 
        .CO(\CARRYB[12][20] ), .S(\SUMB[12][20] ) );
  FA_X1 S2_12_21 ( .A(\CARRYB[11][21] ), .B(\ab[12][21] ), .CI(\SUMB[11][22] ), 
        .CO(\CARRYB[12][21] ), .S(\SUMB[12][21] ) );
  FA_X1 S2_12_22 ( .A(\ab[12][22] ), .B(\CARRYB[11][22] ), .CI(\SUMB[11][23] ), 
        .CO(\CARRYB[12][22] ), .S(\SUMB[12][22] ) );
  FA_X1 S2_12_23 ( .A(\ab[12][23] ), .B(\CARRYB[11][23] ), .CI(\SUMB[11][24] ), 
        .CO(\CARRYB[12][23] ), .S(\SUMB[12][23] ) );
  FA_X1 S2_12_24 ( .A(\ab[12][24] ), .B(\CARRYB[11][24] ), .CI(\SUMB[11][25] ), 
        .CO(\CARRYB[12][24] ), .S(\SUMB[12][24] ) );
  FA_X1 S2_12_25 ( .A(\ab[12][25] ), .B(\CARRYB[11][25] ), .CI(\SUMB[11][26] ), 
        .CO(\CARRYB[12][25] ), .S(\SUMB[12][25] ) );
  FA_X1 S2_12_26 ( .A(\ab[12][26] ), .B(\CARRYB[11][26] ), .CI(\SUMB[11][27] ), 
        .CO(\CARRYB[12][26] ), .S(\SUMB[12][26] ) );
  FA_X1 S2_12_27 ( .A(\ab[12][27] ), .B(\CARRYB[11][27] ), .CI(\SUMB[11][28] ), 
        .CO(\CARRYB[12][27] ), .S(\SUMB[12][27] ) );
  FA_X1 S2_12_28 ( .A(\ab[12][28] ), .B(\CARRYB[11][28] ), .CI(\SUMB[11][29] ), 
        .CO(\CARRYB[12][28] ), .S(\SUMB[12][28] ) );
  FA_X1 S2_12_29 ( .A(\ab[12][29] ), .B(\CARRYB[11][29] ), .CI(\SUMB[11][30] ), 
        .CO(\CARRYB[12][29] ), .S(\SUMB[12][29] ) );
  FA_X1 S3_12_30 ( .A(\ab[12][30] ), .B(\CARRYB[11][30] ), .CI(\ab[11][31] ), 
        .CO(\CARRYB[12][30] ), .S(\SUMB[12][30] ) );
  FA_X1 S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FA_X1 S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA_X1 S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA_X1 S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA_X1 S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA_X1 S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA_X1 S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA_X1 S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA_X1 S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA_X1 S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA_X1 S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA_X1 S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA_X1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA_X1 S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA_X1 S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA_X1 S2_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\SUMB[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA_X1 S2_11_16 ( .A(\ab[11][16] ), .B(\CARRYB[10][16] ), .CI(\SUMB[10][17] ), 
        .CO(\CARRYB[11][16] ), .S(\SUMB[11][16] ) );
  FA_X1 S2_11_17 ( .A(\ab[11][17] ), .B(\CARRYB[10][17] ), .CI(\SUMB[10][18] ), 
        .CO(\CARRYB[11][17] ), .S(\SUMB[11][17] ) );
  FA_X1 S2_11_18 ( .A(\ab[11][18] ), .B(\CARRYB[10][18] ), .CI(\SUMB[10][19] ), 
        .CO(\CARRYB[11][18] ), .S(\SUMB[11][18] ) );
  FA_X1 S2_11_19 ( .A(\ab[11][19] ), .B(\CARRYB[10][19] ), .CI(\SUMB[10][20] ), 
        .CO(\CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FA_X1 S2_11_20 ( .A(\ab[11][20] ), .B(\CARRYB[10][20] ), .CI(\SUMB[10][21] ), 
        .CO(\CARRYB[11][20] ), .S(\SUMB[11][20] ) );
  FA_X1 S2_11_21 ( .A(\ab[11][21] ), .B(\CARRYB[10][21] ), .CI(\SUMB[10][22] ), 
        .CO(\CARRYB[11][21] ), .S(\SUMB[11][21] ) );
  FA_X1 S2_11_22 ( .A(\ab[11][22] ), .B(\CARRYB[10][22] ), .CI(\SUMB[10][23] ), 
        .CO(\CARRYB[11][22] ), .S(\SUMB[11][22] ) );
  FA_X1 S2_11_23 ( .A(\CARRYB[10][23] ), .B(\ab[11][23] ), .CI(\SUMB[10][24] ), 
        .CO(\CARRYB[11][23] ), .S(\SUMB[11][23] ) );
  FA_X1 S2_11_24 ( .A(\ab[11][24] ), .B(\CARRYB[10][24] ), .CI(\SUMB[10][25] ), 
        .CO(\CARRYB[11][24] ), .S(\SUMB[11][24] ) );
  FA_X1 S2_11_25 ( .A(\ab[11][25] ), .B(\CARRYB[10][25] ), .CI(\SUMB[10][26] ), 
        .CO(\CARRYB[11][25] ), .S(\SUMB[11][25] ) );
  FA_X1 S2_11_26 ( .A(\ab[11][26] ), .B(\CARRYB[10][26] ), .CI(\SUMB[10][27] ), 
        .CO(\CARRYB[11][26] ), .S(\SUMB[11][26] ) );
  FA_X1 S2_11_27 ( .A(\ab[11][27] ), .B(\CARRYB[10][27] ), .CI(\SUMB[10][28] ), 
        .CO(\CARRYB[11][27] ), .S(\SUMB[11][27] ) );
  FA_X1 S2_11_28 ( .A(\ab[11][28] ), .B(\CARRYB[10][28] ), .CI(\SUMB[10][29] ), 
        .CO(\CARRYB[11][28] ), .S(\SUMB[11][28] ) );
  FA_X1 S2_11_29 ( .A(\ab[11][29] ), .B(\CARRYB[10][29] ), .CI(\SUMB[10][30] ), 
        .CO(\CARRYB[11][29] ), .S(\SUMB[11][29] ) );
  FA_X1 S3_11_30 ( .A(\ab[11][30] ), .B(\CARRYB[10][30] ), .CI(\ab[10][31] ), 
        .CO(\CARRYB[11][30] ), .S(\SUMB[11][30] ) );
  FA_X1 S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA_X1 S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA_X1 S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA_X1 S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA_X1 S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA_X1 S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA_X1 S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA_X1 S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA_X1 S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA_X1 S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA_X1 S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA_X1 S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA_X1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA_X1 S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA_X1 S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA_X1 S2_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(\SUMB[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA_X1 S2_10_16 ( .A(\ab[10][16] ), .B(\CARRYB[9][16] ), .CI(\SUMB[9][17] ), 
        .CO(\CARRYB[10][16] ), .S(\SUMB[10][16] ) );
  FA_X1 S2_10_17 ( .A(\ab[10][17] ), .B(\CARRYB[9][17] ), .CI(\SUMB[9][18] ), 
        .CO(\CARRYB[10][17] ), .S(\SUMB[10][17] ) );
  FA_X1 S2_10_18 ( .A(\ab[10][18] ), .B(\CARRYB[9][18] ), .CI(\SUMB[9][19] ), 
        .CO(\CARRYB[10][18] ), .S(\SUMB[10][18] ) );
  FA_X1 S2_10_19 ( .A(\ab[10][19] ), .B(\CARRYB[9][19] ), .CI(\SUMB[9][20] ), 
        .CO(\CARRYB[10][19] ), .S(\SUMB[10][19] ) );
  FA_X1 S2_10_20 ( .A(\ab[10][20] ), .B(\CARRYB[9][20] ), .CI(\SUMB[9][21] ), 
        .CO(\CARRYB[10][20] ), .S(\SUMB[10][20] ) );
  FA_X1 S2_10_21 ( .A(\ab[10][21] ), .B(\CARRYB[9][21] ), .CI(\SUMB[9][22] ), 
        .CO(\CARRYB[10][21] ), .S(\SUMB[10][21] ) );
  FA_X1 S2_10_22 ( .A(\ab[10][22] ), .B(\CARRYB[9][22] ), .CI(\SUMB[9][23] ), 
        .CO(\CARRYB[10][22] ), .S(\SUMB[10][22] ) );
  FA_X1 S2_10_23 ( .A(\CARRYB[9][23] ), .B(\ab[10][23] ), .CI(\SUMB[9][24] ), 
        .CO(\CARRYB[10][23] ), .S(\SUMB[10][23] ) );
  FA_X1 S2_10_24 ( .A(\ab[10][24] ), .B(\CARRYB[9][24] ), .CI(\SUMB[9][25] ), 
        .CO(\CARRYB[10][24] ), .S(\SUMB[10][24] ) );
  FA_X1 S2_10_25 ( .A(\ab[10][25] ), .B(\CARRYB[9][25] ), .CI(\SUMB[9][26] ), 
        .CO(\CARRYB[10][25] ), .S(\SUMB[10][25] ) );
  FA_X1 S2_10_26 ( .A(\ab[10][26] ), .B(\CARRYB[9][26] ), .CI(\SUMB[9][27] ), 
        .CO(\CARRYB[10][26] ), .S(\SUMB[10][26] ) );
  FA_X1 S2_10_27 ( .A(\ab[10][27] ), .B(\CARRYB[9][27] ), .CI(\SUMB[9][28] ), 
        .CO(\CARRYB[10][27] ), .S(\SUMB[10][27] ) );
  FA_X1 S2_10_28 ( .A(\ab[10][28] ), .B(\CARRYB[9][28] ), .CI(\SUMB[9][29] ), 
        .CO(\CARRYB[10][28] ), .S(\SUMB[10][28] ) );
  FA_X1 S2_10_29 ( .A(\ab[10][29] ), .B(\CARRYB[9][29] ), .CI(\SUMB[9][30] ), 
        .CO(\CARRYB[10][29] ), .S(\SUMB[10][29] ) );
  FA_X1 S3_10_30 ( .A(\ab[10][30] ), .B(\CARRYB[9][30] ), .CI(\ab[9][31] ), 
        .CO(\CARRYB[10][30] ), .S(\SUMB[10][30] ) );
  FA_X1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA_X1 S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA_X1 S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA_X1 S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA_X1 S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA_X1 S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA_X1 S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA_X1 S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA_X1 S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA_X1 S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA_X1 S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA_X1 S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA_X1 S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA_X1 S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA_X1 S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA_X1 S2_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\SUMB[8][16] ), 
        .CO(\CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA_X1 S2_9_16 ( .A(\ab[9][16] ), .B(\CARRYB[8][16] ), .CI(\SUMB[8][17] ), 
        .CO(\CARRYB[9][16] ), .S(\SUMB[9][16] ) );
  FA_X1 S2_9_17 ( .A(\ab[9][17] ), .B(\CARRYB[8][17] ), .CI(\SUMB[8][18] ), 
        .CO(\CARRYB[9][17] ), .S(\SUMB[9][17] ) );
  FA_X1 S2_9_18 ( .A(\ab[9][18] ), .B(\CARRYB[8][18] ), .CI(\SUMB[8][19] ), 
        .CO(\CARRYB[9][18] ), .S(\SUMB[9][18] ) );
  FA_X1 S2_9_19 ( .A(\ab[9][19] ), .B(\CARRYB[8][19] ), .CI(\SUMB[8][20] ), 
        .CO(\CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FA_X1 S2_9_20 ( .A(\ab[9][20] ), .B(\CARRYB[8][20] ), .CI(\SUMB[8][21] ), 
        .CO(\CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FA_X1 S2_9_21 ( .A(\ab[9][21] ), .B(\CARRYB[8][21] ), .CI(\SUMB[8][22] ), 
        .CO(\CARRYB[9][21] ), .S(\SUMB[9][21] ) );
  FA_X1 S2_9_22 ( .A(\ab[9][22] ), .B(\CARRYB[8][22] ), .CI(\SUMB[8][23] ), 
        .CO(\CARRYB[9][22] ), .S(\SUMB[9][22] ) );
  FA_X1 S2_9_23 ( .A(\CARRYB[8][23] ), .B(\ab[9][23] ), .CI(\SUMB[8][24] ), 
        .CO(\CARRYB[9][23] ), .S(\SUMB[9][23] ) );
  FA_X1 S2_9_24 ( .A(\ab[9][24] ), .B(\CARRYB[8][24] ), .CI(\SUMB[8][25] ), 
        .CO(\CARRYB[9][24] ), .S(\SUMB[9][24] ) );
  FA_X1 S2_9_25 ( .A(\CARRYB[8][25] ), .B(\ab[9][25] ), .CI(\SUMB[8][26] ), 
        .CO(\CARRYB[9][25] ), .S(\SUMB[9][25] ) );
  FA_X1 S2_9_26 ( .A(\ab[9][26] ), .B(\CARRYB[8][26] ), .CI(\SUMB[8][27] ), 
        .CO(\CARRYB[9][26] ), .S(\SUMB[9][26] ) );
  FA_X1 S2_9_27 ( .A(\ab[9][27] ), .B(\CARRYB[8][27] ), .CI(\SUMB[8][28] ), 
        .CO(\CARRYB[9][27] ), .S(\SUMB[9][27] ) );
  FA_X1 S2_9_28 ( .A(\ab[9][28] ), .B(\CARRYB[8][28] ), .CI(\SUMB[8][29] ), 
        .CO(\CARRYB[9][28] ), .S(\SUMB[9][28] ) );
  FA_X1 S2_9_29 ( .A(\ab[9][29] ), .B(\CARRYB[8][29] ), .CI(\SUMB[8][30] ), 
        .CO(\CARRYB[9][29] ), .S(\SUMB[9][29] ) );
  FA_X1 S3_9_30 ( .A(\ab[9][30] ), .B(\CARRYB[8][30] ), .CI(\ab[8][31] ), .CO(
        \CARRYB[9][30] ), .S(\SUMB[9][30] ) );
  FA_X1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA_X1 S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA_X1 S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA_X1 S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA_X1 S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA_X1 S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA_X1 S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA_X1 S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA_X1 S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA_X1 S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA_X1 S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA_X1 S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA_X1 S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA_X1 S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA_X1 S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA_X1 S2_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), 
        .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA_X1 S2_8_16 ( .A(\ab[8][16] ), .B(\CARRYB[7][16] ), .CI(\SUMB[7][17] ), 
        .CO(\CARRYB[8][16] ), .S(\SUMB[8][16] ) );
  FA_X1 S2_8_17 ( .A(\ab[8][17] ), .B(\CARRYB[7][17] ), .CI(\SUMB[7][18] ), 
        .CO(\CARRYB[8][17] ), .S(\SUMB[8][17] ) );
  FA_X1 S2_8_18 ( .A(\ab[8][18] ), .B(\CARRYB[7][18] ), .CI(\SUMB[7][19] ), 
        .CO(\CARRYB[8][18] ), .S(\SUMB[8][18] ) );
  FA_X1 S2_8_19 ( .A(\ab[8][19] ), .B(\CARRYB[7][19] ), .CI(\SUMB[7][20] ), 
        .CO(\CARRYB[8][19] ), .S(\SUMB[8][19] ) );
  FA_X1 S2_8_20 ( .A(\ab[8][20] ), .B(\CARRYB[7][20] ), .CI(\SUMB[7][21] ), 
        .CO(\CARRYB[8][20] ), .S(\SUMB[8][20] ) );
  FA_X1 S2_8_21 ( .A(\ab[8][21] ), .B(\CARRYB[7][21] ), .CI(\SUMB[7][22] ), 
        .CO(\CARRYB[8][21] ), .S(\SUMB[8][21] ) );
  FA_X1 S2_8_22 ( .A(\ab[8][22] ), .B(\CARRYB[7][22] ), .CI(\SUMB[7][23] ), 
        .CO(\CARRYB[8][22] ), .S(\SUMB[8][22] ) );
  FA_X1 S2_8_23 ( .A(\ab[8][23] ), .B(\CARRYB[7][23] ), .CI(\SUMB[7][24] ), 
        .CO(\CARRYB[8][23] ), .S(\SUMB[8][23] ) );
  FA_X1 S2_8_24 ( .A(\ab[8][24] ), .B(\CARRYB[7][24] ), .CI(\SUMB[7][25] ), 
        .CO(\CARRYB[8][24] ), .S(\SUMB[8][24] ) );
  FA_X1 S2_8_25 ( .A(\ab[8][25] ), .B(\CARRYB[7][25] ), .CI(\SUMB[7][26] ), 
        .CO(\CARRYB[8][25] ), .S(\SUMB[8][25] ) );
  FA_X1 S2_8_26 ( .A(\ab[8][26] ), .B(\CARRYB[7][26] ), .CI(\SUMB[7][27] ), 
        .CO(\CARRYB[8][26] ), .S(\SUMB[8][26] ) );
  FA_X1 S2_8_27 ( .A(\ab[8][27] ), .B(\CARRYB[7][27] ), .CI(\SUMB[7][28] ), 
        .CO(\CARRYB[8][27] ), .S(\SUMB[8][27] ) );
  FA_X1 S2_8_28 ( .A(\ab[8][28] ), .B(\CARRYB[7][28] ), .CI(\SUMB[7][29] ), 
        .CO(\CARRYB[8][28] ), .S(\SUMB[8][28] ) );
  FA_X1 S2_8_29 ( .A(\ab[8][29] ), .B(\CARRYB[7][29] ), .CI(\SUMB[7][30] ), 
        .CO(\CARRYB[8][29] ), .S(\SUMB[8][29] ) );
  FA_X1 S3_8_30 ( .A(\ab[8][30] ), .B(\CARRYB[7][30] ), .CI(\ab[7][31] ), .CO(
        \CARRYB[8][30] ), .S(\SUMB[8][30] ) );
  FA_X1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA_X1 S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA_X1 S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA_X1 S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA_X1 S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA_X1 S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA_X1 S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA_X1 S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA_X1 S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA_X1 S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA_X1 S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA_X1 S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA_X1 S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA_X1 S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA_X1 S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA_X1 S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), 
        .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA_X1 S2_7_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .CI(\SUMB[6][17] ), 
        .CO(\CARRYB[7][16] ), .S(\SUMB[7][16] ) );
  FA_X1 S2_7_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .CI(\SUMB[6][18] ), 
        .CO(\CARRYB[7][17] ), .S(\SUMB[7][17] ) );
  FA_X1 S2_7_18 ( .A(\CARRYB[6][18] ), .B(\ab[7][18] ), .CI(\SUMB[6][19] ), 
        .CO(\CARRYB[7][18] ), .S(\SUMB[7][18] ) );
  FA_X1 S2_7_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .CI(\SUMB[6][20] ), 
        .CO(\CARRYB[7][19] ), .S(\SUMB[7][19] ) );
  FA_X1 S2_7_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .CI(\SUMB[6][21] ), 
        .CO(\CARRYB[7][20] ), .S(\SUMB[7][20] ) );
  FA_X1 S2_7_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .CI(\SUMB[6][22] ), 
        .CO(\CARRYB[7][21] ), .S(\SUMB[7][21] ) );
  FA_X1 S2_7_22 ( .A(\ab[7][22] ), .B(\CARRYB[6][22] ), .CI(\SUMB[6][23] ), 
        .CO(\CARRYB[7][22] ), .S(\SUMB[7][22] ) );
  FA_X1 S2_7_23 ( .A(\ab[7][23] ), .B(\CARRYB[6][23] ), .CI(\SUMB[6][24] ), 
        .CO(\CARRYB[7][23] ), .S(\SUMB[7][23] ) );
  FA_X1 S2_7_24 ( .A(\ab[7][24] ), .B(\CARRYB[6][24] ), .CI(\SUMB[6][25] ), 
        .CO(\CARRYB[7][24] ), .S(\SUMB[7][24] ) );
  FA_X1 S2_7_25 ( .A(\ab[7][25] ), .B(\CARRYB[6][25] ), .CI(\SUMB[6][26] ), 
        .CO(\CARRYB[7][25] ), .S(\SUMB[7][25] ) );
  FA_X1 S2_7_26 ( .A(\ab[7][26] ), .B(\CARRYB[6][26] ), .CI(\SUMB[6][27] ), 
        .CO(\CARRYB[7][26] ), .S(\SUMB[7][26] ) );
  FA_X1 S2_7_27 ( .A(\CARRYB[6][27] ), .B(\ab[7][27] ), .CI(\SUMB[6][28] ), 
        .CO(\CARRYB[7][27] ), .S(\SUMB[7][27] ) );
  FA_X1 S2_7_28 ( .A(\ab[7][28] ), .B(\CARRYB[6][28] ), .CI(\SUMB[6][29] ), 
        .CO(\CARRYB[7][28] ), .S(\SUMB[7][28] ) );
  FA_X1 S2_7_29 ( .A(\ab[7][29] ), .B(\CARRYB[6][29] ), .CI(\SUMB[6][30] ), 
        .CO(\CARRYB[7][29] ), .S(\SUMB[7][29] ) );
  FA_X1 S3_7_30 ( .A(\ab[7][30] ), .B(\CARRYB[6][30] ), .CI(\ab[6][31] ), .CO(
        \CARRYB[7][30] ), .S(\SUMB[7][30] ) );
  FA_X1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA_X1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA_X1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA_X1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA_X1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA_X1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA_X1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA_X1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA_X1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA_X1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA_X1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA_X1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA_X1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA_X1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA_X1 S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA_X1 S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\SUMB[5][16] ), 
        .CO(\CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA_X1 S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .CI(\SUMB[5][17] ), 
        .CO(\CARRYB[6][16] ), .S(\SUMB[6][16] ) );
  FA_X1 S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .CI(\SUMB[5][18] ), 
        .CO(\CARRYB[6][17] ), .S(\SUMB[6][17] ) );
  FA_X1 S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .CI(\SUMB[5][19] ), 
        .CO(\CARRYB[6][18] ), .S(\SUMB[6][18] ) );
  FA_X1 S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .CI(\SUMB[5][20] ), 
        .CO(\CARRYB[6][19] ), .S(\SUMB[6][19] ) );
  FA_X1 S2_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .CI(\SUMB[5][21] ), 
        .CO(\CARRYB[6][20] ), .S(\SUMB[6][20] ) );
  FA_X1 S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .CI(\SUMB[5][22] ), 
        .CO(\CARRYB[6][21] ), .S(\SUMB[6][21] ) );
  FA_X1 S2_6_22 ( .A(\ab[6][22] ), .B(\CARRYB[5][22] ), .CI(\SUMB[5][23] ), 
        .CO(\CARRYB[6][22] ), .S(\SUMB[6][22] ) );
  FA_X1 S2_6_23 ( .A(\ab[6][23] ), .B(\CARRYB[5][23] ), .CI(\SUMB[5][24] ), 
        .CO(\CARRYB[6][23] ), .S(\SUMB[6][23] ) );
  FA_X1 S2_6_24 ( .A(\ab[6][24] ), .B(\CARRYB[5][24] ), .CI(\SUMB[5][25] ), 
        .CO(\CARRYB[6][24] ), .S(\SUMB[6][24] ) );
  FA_X1 S2_6_25 ( .A(\ab[6][25] ), .B(\CARRYB[5][25] ), .CI(\SUMB[5][26] ), 
        .CO(\CARRYB[6][25] ), .S(\SUMB[6][25] ) );
  FA_X1 S2_6_26 ( .A(\ab[6][26] ), .B(\CARRYB[5][26] ), .CI(\SUMB[5][27] ), 
        .CO(\CARRYB[6][26] ), .S(\SUMB[6][26] ) );
  FA_X1 S2_6_27 ( .A(\ab[6][27] ), .B(\CARRYB[5][27] ), .CI(\SUMB[5][28] ), 
        .CO(\CARRYB[6][27] ), .S(\SUMB[6][27] ) );
  FA_X1 S2_6_28 ( .A(\ab[6][28] ), .B(\CARRYB[5][28] ), .CI(\SUMB[5][29] ), 
        .CO(\CARRYB[6][28] ), .S(\SUMB[6][28] ) );
  FA_X1 S2_6_29 ( .A(\ab[6][29] ), .B(\CARRYB[5][29] ), .CI(\SUMB[5][30] ), 
        .CO(\CARRYB[6][29] ), .S(\SUMB[6][29] ) );
  FA_X1 S3_6_30 ( .A(\ab[6][30] ), .B(\CARRYB[5][30] ), .CI(\ab[5][31] ), .CO(
        \CARRYB[6][30] ), .S(\SUMB[6][30] ) );
  FA_X1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA_X1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA_X1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA_X1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA_X1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA_X1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA_X1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA_X1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA_X1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA_X1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA_X1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA_X1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA_X1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA_X1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA_X1 S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA_X1 S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), 
        .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA_X1 S2_5_16 ( .A(\ab[5][16] ), .B(\CARRYB[4][16] ), .CI(\SUMB[4][17] ), 
        .CO(\CARRYB[5][16] ), .S(\SUMB[5][16] ) );
  FA_X1 S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .CI(\SUMB[4][18] ), 
        .CO(\CARRYB[5][17] ), .S(\SUMB[5][17] ) );
  FA_X1 S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .CI(\SUMB[4][19] ), 
        .CO(\CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FA_X1 S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .CI(\SUMB[4][20] ), 
        .CO(\CARRYB[5][19] ), .S(\SUMB[5][19] ) );
  FA_X1 S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .CI(\SUMB[4][21] ), 
        .CO(\CARRYB[5][20] ), .S(\SUMB[5][20] ) );
  FA_X1 S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .CI(\SUMB[4][22] ), 
        .CO(\CARRYB[5][21] ), .S(\SUMB[5][21] ) );
  FA_X1 S2_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .CI(\SUMB[4][23] ), 
        .CO(\CARRYB[5][22] ), .S(\SUMB[5][22] ) );
  FA_X1 S2_5_23 ( .A(\ab[5][23] ), .B(\CARRYB[4][23] ), .CI(\SUMB[4][24] ), 
        .CO(\CARRYB[5][23] ), .S(\SUMB[5][23] ) );
  FA_X1 S2_5_24 ( .A(\ab[5][24] ), .B(\CARRYB[4][24] ), .CI(\SUMB[4][25] ), 
        .CO(\CARRYB[5][24] ), .S(\SUMB[5][24] ) );
  FA_X1 S2_5_25 ( .A(\ab[5][25] ), .B(\CARRYB[4][25] ), .CI(\SUMB[4][26] ), 
        .CO(\CARRYB[5][25] ), .S(\SUMB[5][25] ) );
  FA_X1 S2_5_26 ( .A(\ab[5][26] ), .B(\CARRYB[4][26] ), .CI(\SUMB[4][27] ), 
        .CO(\CARRYB[5][26] ), .S(\SUMB[5][26] ) );
  FA_X1 S2_5_27 ( .A(\ab[5][27] ), .B(\CARRYB[4][27] ), .CI(\SUMB[4][28] ), 
        .CO(\CARRYB[5][27] ), .S(\SUMB[5][27] ) );
  FA_X1 S2_5_28 ( .A(\ab[5][28] ), .B(\CARRYB[4][28] ), .CI(\SUMB[4][29] ), 
        .CO(\CARRYB[5][28] ), .S(\SUMB[5][28] ) );
  FA_X1 S2_5_29 ( .A(\CARRYB[4][29] ), .B(\ab[5][29] ), .CI(\SUMB[4][30] ), 
        .CO(\CARRYB[5][29] ), .S(\SUMB[5][29] ) );
  FA_X1 S3_5_30 ( .A(\ab[5][30] ), .B(\CARRYB[4][30] ), .CI(\ab[4][31] ), .CO(
        \CARRYB[5][30] ), .S(\SUMB[5][30] ) );
  FA_X1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA_X1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA_X1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA_X1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA_X1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA_X1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA_X1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA_X1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA_X1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA_X1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA_X1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA_X1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA_X1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA_X1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA_X1 S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA_X1 S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), 
        .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA_X1 S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .CI(\SUMB[3][17] ), 
        .CO(\CARRYB[4][16] ), .S(\SUMB[4][16] ) );
  FA_X1 S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .CI(\SUMB[3][18] ), 
        .CO(\CARRYB[4][17] ), .S(\SUMB[4][17] ) );
  FA_X1 S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .CI(\SUMB[3][19] ), 
        .CO(\CARRYB[4][18] ), .S(\SUMB[4][18] ) );
  FA_X1 S2_4_19 ( .A(\ab[4][19] ), .B(\CARRYB[3][19] ), .CI(\SUMB[3][20] ), 
        .CO(\CARRYB[4][19] ), .S(\SUMB[4][19] ) );
  FA_X1 S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .CI(\SUMB[3][21] ), 
        .CO(\CARRYB[4][20] ), .S(\SUMB[4][20] ) );
  FA_X1 S2_4_21 ( .A(\ab[4][21] ), .B(\CARRYB[3][21] ), .CI(\SUMB[3][22] ), 
        .CO(\CARRYB[4][21] ), .S(\SUMB[4][21] ) );
  FA_X1 S2_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .CI(\SUMB[3][23] ), 
        .CO(\CARRYB[4][22] ), .S(\SUMB[4][22] ) );
  FA_X1 S2_4_23 ( .A(\ab[4][23] ), .B(\CARRYB[3][23] ), .CI(\SUMB[3][24] ), 
        .CO(\CARRYB[4][23] ), .S(\SUMB[4][23] ) );
  FA_X1 S2_4_24 ( .A(\ab[4][24] ), .B(\CARRYB[3][24] ), .CI(\SUMB[3][25] ), 
        .CO(\CARRYB[4][24] ), .S(\SUMB[4][24] ) );
  FA_X1 S2_4_25 ( .A(\ab[4][25] ), .B(\CARRYB[3][25] ), .CI(\SUMB[3][26] ), 
        .CO(\CARRYB[4][25] ), .S(\SUMB[4][25] ) );
  FA_X1 S2_4_26 ( .A(\ab[4][26] ), .B(\CARRYB[3][26] ), .CI(\SUMB[3][27] ), 
        .CO(\CARRYB[4][26] ), .S(\SUMB[4][26] ) );
  FA_X1 S2_4_27 ( .A(\ab[4][27] ), .B(\CARRYB[3][27] ), .CI(\SUMB[3][28] ), 
        .CO(\CARRYB[4][27] ), .S(\SUMB[4][27] ) );
  FA_X1 S2_4_28 ( .A(\ab[4][28] ), .B(\CARRYB[3][28] ), .CI(\SUMB[3][29] ), 
        .CO(\CARRYB[4][28] ), .S(\SUMB[4][28] ) );
  FA_X1 S2_4_29 ( .A(\CARRYB[3][29] ), .B(\ab[4][29] ), .CI(\SUMB[3][30] ), 
        .CO(\CARRYB[4][29] ), .S(\SUMB[4][29] ) );
  FA_X1 S3_4_30 ( .A(\ab[4][30] ), .B(\CARRYB[3][30] ), .CI(\ab[3][31] ), .CO(
        \CARRYB[4][30] ), .S(\SUMB[4][30] ) );
  FA_X1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA_X1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA_X1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA_X1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA_X1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA_X1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA_X1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA_X1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA_X1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA_X1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA_X1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA_X1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA_X1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA_X1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA_X1 S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA_X1 S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), 
        .CO(\CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA_X1 S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .CI(\SUMB[2][17] ), 
        .CO(\CARRYB[3][16] ), .S(\SUMB[3][16] ) );
  FA_X1 S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .CI(\SUMB[2][18] ), 
        .CO(\CARRYB[3][17] ), .S(\SUMB[3][17] ) );
  FA_X1 S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .CI(\SUMB[2][19] ), 
        .CO(\CARRYB[3][18] ), .S(\SUMB[3][18] ) );
  FA_X1 S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .CI(\SUMB[2][20] ), 
        .CO(\CARRYB[3][19] ), .S(\SUMB[3][19] ) );
  FA_X1 S2_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .CI(\SUMB[2][21] ), 
        .CO(\CARRYB[3][20] ), .S(\SUMB[3][20] ) );
  FA_X1 S2_3_21 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .CI(\SUMB[2][22] ), 
        .CO(\CARRYB[3][21] ), .S(\SUMB[3][21] ) );
  FA_X1 S2_3_22 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .CI(\SUMB[2][23] ), 
        .CO(\CARRYB[3][22] ), .S(\SUMB[3][22] ) );
  FA_X1 S2_3_23 ( .A(\ab[3][23] ), .B(\CARRYB[2][23] ), .CI(\SUMB[2][24] ), 
        .CO(\CARRYB[3][23] ), .S(\SUMB[3][23] ) );
  FA_X1 S2_3_24 ( .A(\ab[3][24] ), .B(\CARRYB[2][24] ), .CI(\SUMB[2][25] ), 
        .CO(\CARRYB[3][24] ), .S(\SUMB[3][24] ) );
  FA_X1 S2_3_25 ( .A(\ab[3][25] ), .B(\CARRYB[2][25] ), .CI(\SUMB[2][26] ), 
        .CO(\CARRYB[3][25] ), .S(\SUMB[3][25] ) );
  FA_X1 S2_3_26 ( .A(\ab[3][26] ), .B(\CARRYB[2][26] ), .CI(\SUMB[2][27] ), 
        .CO(\CARRYB[3][26] ), .S(\SUMB[3][26] ) );
  FA_X1 S2_3_27 ( .A(\ab[3][27] ), .B(\CARRYB[2][27] ), .CI(\SUMB[2][28] ), 
        .CO(\CARRYB[3][27] ), .S(\SUMB[3][27] ) );
  FA_X1 S2_3_28 ( .A(\ab[3][28] ), .B(\CARRYB[2][28] ), .CI(\SUMB[2][29] ), 
        .CO(\CARRYB[3][28] ), .S(\SUMB[3][28] ) );
  FA_X1 S2_3_29 ( .A(\CARRYB[2][29] ), .B(\ab[3][29] ), .CI(\SUMB[2][30] ), 
        .CO(\CARRYB[3][29] ), .S(\SUMB[3][29] ) );
  FA_X1 S3_3_30 ( .A(\ab[3][30] ), .B(\CARRYB[2][30] ), .CI(\ab[2][31] ), .CO(
        \CARRYB[3][30] ), .S(\SUMB[3][30] ) );
  FA_X1 S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA_X1 S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA_X1 S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA_X1 S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA_X1 S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA_X1 S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA_X1 S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA_X1 S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA_X1 S2_2_10 ( .A(\ab[2][10] ), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), 
        .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FA_X1 S2_2_11 ( .A(\ab[2][11] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), 
        .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FA_X1 S2_2_12 ( .A(\ab[2][12] ), .B(\CARRYB[1][12] ), .CI(\SUMB[1][13] ), 
        .CO(\CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FA_X1 S2_2_13 ( .A(\ab[2][13] ), .B(\CARRYB[1][13] ), .CI(\SUMB[1][14] ), 
        .CO(\CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FA_X1 S2_2_14 ( .A(\ab[2][14] ), .B(\CARRYB[1][14] ), .CI(\SUMB[1][15] ), 
        .CO(\CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  FA_X1 S2_2_15 ( .A(\ab[2][15] ), .B(\CARRYB[1][15] ), .CI(\SUMB[1][16] ), 
        .CO(\CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  FA_X1 S2_2_16 ( .A(\ab[2][16] ), .B(\CARRYB[1][16] ), .CI(\SUMB[1][17] ), 
        .CO(\CARRYB[2][16] ), .S(\SUMB[2][16] ) );
  FA_X1 S2_2_17 ( .A(\ab[2][17] ), .B(\CARRYB[1][17] ), .CI(\SUMB[1][18] ), 
        .CO(\CARRYB[2][17] ), .S(\SUMB[2][17] ) );
  FA_X1 S2_2_18 ( .A(\ab[2][18] ), .B(\CARRYB[1][18] ), .CI(\SUMB[1][19] ), 
        .CO(\CARRYB[2][18] ), .S(\SUMB[2][18] ) );
  FA_X1 S2_2_19 ( .A(\ab[2][19] ), .B(\CARRYB[1][19] ), .CI(\SUMB[1][20] ), 
        .CO(\CARRYB[2][19] ), .S(\SUMB[2][19] ) );
  FA_X1 S2_2_20 ( .A(\ab[2][20] ), .B(\CARRYB[1][20] ), .CI(\SUMB[1][21] ), 
        .CO(\CARRYB[2][20] ), .S(\SUMB[2][20] ) );
  FA_X1 S2_2_21 ( .A(\ab[2][21] ), .B(\CARRYB[1][21] ), .CI(\SUMB[1][22] ), 
        .CO(\CARRYB[2][21] ), .S(\SUMB[2][21] ) );
  FA_X1 S2_2_22 ( .A(\ab[2][22] ), .B(\CARRYB[1][22] ), .CI(\SUMB[1][23] ), 
        .CO(\CARRYB[2][22] ), .S(\SUMB[2][22] ) );
  FA_X1 S2_2_23 ( .A(\ab[2][23] ), .B(\CARRYB[1][23] ), .CI(\SUMB[1][24] ), 
        .CO(\CARRYB[2][23] ), .S(\SUMB[2][23] ) );
  FA_X1 S2_2_24 ( .A(\ab[2][24] ), .B(\CARRYB[1][24] ), .CI(\SUMB[1][25] ), 
        .CO(\CARRYB[2][24] ), .S(\SUMB[2][24] ) );
  FA_X1 S2_2_25 ( .A(\SUMB[1][26] ), .B(\CARRYB[1][25] ), .CI(\ab[2][25] ), 
        .CO(\CARRYB[2][25] ), .S(\SUMB[2][25] ) );
  FA_X1 S2_2_26 ( .A(\ab[2][26] ), .B(\CARRYB[1][26] ), .CI(\SUMB[1][27] ), 
        .CO(\CARRYB[2][26] ), .S(\SUMB[2][26] ) );
  FA_X1 S2_2_27 ( .A(\CARRYB[1][27] ), .B(\ab[2][27] ), .CI(\SUMB[1][28] ), 
        .CO(\CARRYB[2][27] ), .S(\SUMB[2][27] ) );
  FA_X1 S2_2_28 ( .A(\SUMB[1][29] ), .B(\CARRYB[1][28] ), .CI(\ab[2][28] ), 
        .CO(\CARRYB[2][28] ), .S(\SUMB[2][28] ) );
  FA_X1 S2_2_29 ( .A(\ab[2][29] ), .B(\CARRYB[1][29] ), .CI(\SUMB[1][30] ), 
        .CO(\CARRYB[2][29] ), .S(\SUMB[2][29] ) );
  FA_X1 S3_2_30 ( .A(\ab[1][31] ), .B(\CARRYB[1][30] ), .CI(\ab[2][30] ), .CO(
        \CARRYB[2][30] ), .S(\SUMB[2][30] ) );
  XOR2_X1 U67 ( .A(\CARRYB[31][10] ), .B(\SUMB[31][11] ), .Z(\A1[40] ) );
  XOR2_X1 U69 ( .A(\CARRYB[31][11] ), .B(\SUMB[31][12] ), .Z(\A1[41] ) );
  XOR2_X1 U71 ( .A(\CARRYB[31][13] ), .B(\SUMB[31][14] ), .Z(\A1[43] ) );
  XOR2_X1 U73 ( .A(\CARRYB[31][12] ), .B(\SUMB[31][13] ), .Z(\A1[42] ) );
  XOR2_X1 U75 ( .A(\SUMB[31][1] ), .B(\CARRYB[31][0] ), .Z(\A1[30] ) );
  XOR2_X1 U77 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Z(PRODUCT[1]) );
  XOR2_X1 U79 ( .A(\CARRYB[31][1] ), .B(\SUMB[31][2] ), .Z(\A1[31] ) );
  XOR2_X1 U81 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(\SUMB[1][1] ) );
  XOR2_X1 U83 ( .A(\SUMB[31][4] ), .B(\CARRYB[31][3] ), .Z(\A1[33] ) );
  XOR2_X1 U87 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(\SUMB[1][3] ) );
  XOR2_X1 U89 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(\SUMB[1][2] ) );
  XOR2_X1 U91 ( .A(\CARRYB[31][4] ), .B(\SUMB[31][5] ), .Z(\A1[34] ) );
  XOR2_X1 U93 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(\SUMB[1][4] ) );
  XOR2_X1 U95 ( .A(\CARRYB[31][5] ), .B(\SUMB[31][6] ), .Z(\A1[35] ) );
  XOR2_X1 U97 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(\SUMB[1][5] ) );
  XOR2_X1 U99 ( .A(\CARRYB[31][6] ), .B(\SUMB[31][7] ), .Z(\A1[36] ) );
  XOR2_X1 U101 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(\SUMB[1][6] ) );
  XOR2_X1 U103 ( .A(\CARRYB[31][7] ), .B(\SUMB[31][8] ), .Z(\A1[37] ) );
  XOR2_X1 U105 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(\SUMB[1][7] ) );
  XOR2_X1 U107 ( .A(\CARRYB[31][9] ), .B(\SUMB[31][10] ), .Z(\A1[39] ) );
  XOR2_X1 U109 ( .A(\CARRYB[31][8] ), .B(\SUMB[31][9] ), .Z(\A1[38] ) );
  XOR2_X1 U111 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(\SUMB[1][13] ) );
  XOR2_X1 U113 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(\SUMB[1][12] ) );
  XOR2_X1 U115 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(\SUMB[1][11] ) );
  XOR2_X1 U117 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(\SUMB[1][10] ) );
  XOR2_X1 U119 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(\SUMB[1][9] ) );
  XOR2_X1 U121 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(\SUMB[1][8] ) );
  XOR2_X1 U123 ( .A(\CARRYB[31][15] ), .B(\SUMB[31][16] ), .Z(\A1[45] ) );
  XOR2_X1 U125 ( .A(\CARRYB[31][14] ), .B(\SUMB[31][15] ), .Z(\A1[44] ) );
  XOR2_X1 U127 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(\SUMB[1][15] ) );
  XOR2_X1 U129 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(\SUMB[1][14] ) );
  XOR2_X1 U131 ( .A(\CARRYB[31][16] ), .B(\SUMB[31][17] ), .Z(\A1[46] ) );
  XOR2_X1 U133 ( .A(\ab[1][16] ), .B(\ab[0][17] ), .Z(\SUMB[1][16] ) );
  XOR2_X1 U135 ( .A(\CARRYB[31][17] ), .B(\SUMB[31][18] ), .Z(\A1[47] ) );
  XOR2_X1 U137 ( .A(\ab[1][17] ), .B(\ab[0][18] ), .Z(\SUMB[1][17] ) );
  XOR2_X1 U139 ( .A(\CARRYB[31][18] ), .B(\SUMB[31][19] ), .Z(\A1[48] ) );
  XOR2_X1 U141 ( .A(\ab[1][18] ), .B(\ab[0][19] ), .Z(\SUMB[1][18] ) );
  XOR2_X1 U143 ( .A(\CARRYB[31][19] ), .B(\SUMB[31][20] ), .Z(\A1[49] ) );
  XOR2_X1 U145 ( .A(\ab[1][19] ), .B(\ab[0][20] ), .Z(\SUMB[1][19] ) );
  XOR2_X1 U147 ( .A(\CARRYB[31][20] ), .B(\SUMB[31][21] ), .Z(\A1[50] ) );
  XOR2_X1 U149 ( .A(\ab[1][20] ), .B(\ab[0][21] ), .Z(\SUMB[1][20] ) );
  XOR2_X1 U151 ( .A(\CARRYB[31][21] ), .B(\SUMB[31][22] ), .Z(\A1[51] ) );
  XOR2_X1 U153 ( .A(\ab[1][21] ), .B(\ab[0][22] ), .Z(\SUMB[1][21] ) );
  XOR2_X1 U155 ( .A(\CARRYB[31][22] ), .B(\SUMB[31][23] ), .Z(\A1[52] ) );
  XOR2_X1 U159 ( .A(\CARRYB[31][23] ), .B(\SUMB[31][24] ), .Z(\A1[53] ) );
  XOR2_X1 U163 ( .A(\CARRYB[31][24] ), .B(\SUMB[31][25] ), .Z(\A1[54] ) );
  XOR2_X1 U165 ( .A(\ab[1][24] ), .B(\ab[0][25] ), .Z(\SUMB[1][24] ) );
  XOR2_X1 U167 ( .A(\CARRYB[31][25] ), .B(\SUMB[31][26] ), .Z(\A1[55] ) );
  XOR2_X1 U169 ( .A(\ab[1][25] ), .B(\ab[0][26] ), .Z(\SUMB[1][25] ) );
  XOR2_X1 U171 ( .A(\CARRYB[31][26] ), .B(\SUMB[31][27] ), .Z(\A1[56] ) );
  XOR2_X1 U173 ( .A(\ab[1][26] ), .B(\ab[0][27] ), .Z(\SUMB[1][26] ) );
  XOR2_X1 U175 ( .A(\CARRYB[31][27] ), .B(\SUMB[31][28] ), .Z(\A1[57] ) );
  XOR2_X1 U179 ( .A(\CARRYB[31][28] ), .B(\SUMB[31][29] ), .Z(\A1[58] ) );
  XOR2_X1 U181 ( .A(\ab[0][29] ), .B(\ab[1][28] ), .Z(\SUMB[1][28] ) );
  XOR2_X1 U183 ( .A(\CARRYB[31][30] ), .B(\SUMB[31][31] ), .Z(\A1[60] ) );
  XOR2_X1 U185 ( .A(\CARRYB[31][29] ), .B(\SUMB[31][30] ), .Z(\A1[59] ) );
  XOR2_X1 U187 ( .A(\ab[1][30] ), .B(\ab[0][31] ), .Z(\SUMB[1][30] ) );
  Multiplier_NBIT_DATA32_DW01_add_1 FS_1 ( .A({\A1[61] , \A1[60] , \A1[59] , 
        \A1[58] , \A1[57] , \A1[56] , \A1[55] , \A1[54] , \A1[53] , \A1[52] , 
        \A1[51] , \A1[50] , \A1[49] , \A1[48] , \A1[47] , \A1[46] , \A1[45] , 
        \A1[44] , \A1[43] , \A1[42] , \A1[41] , \A1[40] , \A1[39] , \A1[38] , 
        \A1[37] , \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , 
        \A1[30] , \A1[29] , \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , 
        \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , 
        \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , 
        \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , 
        \A1[1] , \A1[0] }), .B({\A2[61] , \A2[60] , \A2[59] , \A2[58] , 
        \A2[57] , \A2[56] , \A2[55] , \A2[54] , \A2[53] , \A2[52] , \A2[51] , 
        \A2[50] , \A2[49] , \A2[48] , \A2[47] , \A2[46] , \A2[45] , \A2[44] , 
        \A2[43] , \A2[42] , \A2[41] , \A2[40] , \A2[39] , \A2[38] , \A2[37] , 
        \A2[36] , \A2[35] , \A2[34] , \A2[33] , \A2[32] , \A2[31] , \A2[30] , 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(PRODUCT[63:2])
         );
  INV_X4 U2 ( .A(A[15]), .ZN(n57) );
  CLKBUF_X3 U3 ( .A(n38), .Z(n110) );
  BUF_X4 U4 ( .A(n8), .Z(n189) );
  CLKBUF_X3 U5 ( .A(n2), .Z(n207) );
  INV_X2 U6 ( .A(A[20]), .ZN(n51) );
  INV_X4 U7 ( .A(A[13]), .ZN(n59) );
  INV_X2 U8 ( .A(A[24]), .ZN(n47) );
  CLKBUF_X3 U9 ( .A(n37), .Z(n112) );
  INV_X2 U10 ( .A(A[23]), .ZN(n48) );
  INV_X2 U11 ( .A(A[22]), .ZN(n49) );
  INV_X2 U12 ( .A(A[18]), .ZN(n54) );
  CLKBUF_X1 U13 ( .A(n16), .Z(n172) );
  BUF_X4 U14 ( .A(n16), .Z(n170) );
  INV_X2 U15 ( .A(A[25]), .ZN(n46) );
  INV_X2 U16 ( .A(A[29]), .ZN(n42) );
  BUF_X4 U17 ( .A(n12), .Z(n180) );
  CLKBUF_X3 U18 ( .A(n36), .Z(n114) );
  INV_X2 U19 ( .A(A[14]), .ZN(n58) );
  CLKBUF_X1 U20 ( .A(n58), .Z(n99) );
  INV_X2 U21 ( .A(A[30]), .ZN(n40) );
  INV_X4 U22 ( .A(A[16]), .ZN(n56) );
  INV_X2 U23 ( .A(A[19]), .ZN(n53) );
  INV_X2 U24 ( .A(A[21]), .ZN(n50) );
  INV_X2 U25 ( .A(A[11]), .ZN(n61) );
  CLKBUF_X3 U26 ( .A(n61), .Z(n97) );
  INV_X2 U27 ( .A(A[28]), .ZN(n43) );
  BUF_X4 U28 ( .A(n62), .Z(n96) );
  INV_X2 U29 ( .A(A[10]), .ZN(n62) );
  BUF_X4 U30 ( .A(n14), .Z(n176) );
  INV_X2 U31 ( .A(A[27]), .ZN(n44) );
  INV_X2 U32 ( .A(A[12]), .ZN(n60) );
  CLKBUF_X3 U33 ( .A(n60), .Z(n98) );
  INV_X2 U34 ( .A(A[26]), .ZN(n45) );
  INV_X2 U35 ( .A(A[17]), .ZN(n55) );
  AND2_X1 U36 ( .A1(n66), .A2(A[2]), .ZN(\ab[2][30] ) );
  CLKBUF_X2 U37 ( .A(n21), .Z(n158) );
  CLKBUF_X3 U38 ( .A(n19), .Z(n164) );
  BUF_X1 U39 ( .A(n63), .Z(n93) );
  BUF_X1 U40 ( .A(n41), .Z(n103) );
  BUF_X1 U41 ( .A(n17), .Z(n168) );
  BUF_X2 U42 ( .A(n5), .Z(n198) );
  CLKBUF_X1 U43 ( .A(B[30]), .Z(n66) );
  BUF_X1 U44 ( .A(n18), .Z(n166) );
  CLKBUF_X1 U45 ( .A(\SUMB[31][4] ), .Z(n67) );
  INV_X1 U46 ( .A(n180), .ZN(n68) );
  NAND2_X1 U47 ( .A1(\ab[1][22] ), .A2(n70), .ZN(n71) );
  NAND2_X1 U48 ( .A1(n69), .A2(\ab[0][23] ), .ZN(n72) );
  NAND2_X1 U49 ( .A1(n71), .A2(n72), .ZN(\SUMB[1][22] ) );
  INV_X1 U50 ( .A(\ab[1][22] ), .ZN(n69) );
  INV_X1 U51 ( .A(\ab[0][23] ), .ZN(n70) );
  CLKBUF_X1 U52 ( .A(n18), .Z(n73) );
  BUF_X1 U53 ( .A(n13), .Z(n178) );
  CLKBUF_X3 U54 ( .A(n20), .Z(n161) );
  CLKBUF_X3 U55 ( .A(n10), .Z(n185) );
  CLKBUF_X1 U56 ( .A(n52), .Z(n100) );
  BUF_X2 U57 ( .A(n92), .Z(n101) );
  CLKBUF_X1 U58 ( .A(n102), .Z(n74) );
  BUF_X2 U59 ( .A(n52), .Z(n102) );
  AND2_X1 U60 ( .A1(B[26]), .A2(n84), .ZN(\ab[0][26] ) );
  BUF_X1 U61 ( .A(A[0]), .Z(n84) );
  XNOR2_X1 U62 ( .A(n75), .B(\ab[0][24] ), .ZN(\SUMB[1][23] ) );
  OR2_X1 U63 ( .A1(n166), .A2(n102), .ZN(n75) );
  NAND2_X1 U64 ( .A1(\ab[1][29] ), .A2(n77), .ZN(n78) );
  NAND2_X1 U65 ( .A1(n76), .A2(\ab[0][30] ), .ZN(n79) );
  NAND2_X1 U66 ( .A1(n78), .A2(n79), .ZN(\SUMB[1][29] ) );
  INV_X1 U68 ( .A(\ab[1][29] ), .ZN(n76) );
  INV_X1 U70 ( .A(\ab[0][30] ), .ZN(n77) );
  CLKBUF_X3 U72 ( .A(n63), .Z(n95) );
  NOR2_X1 U74 ( .A1(n80), .A2(n13), .ZN(\CARRYB[1][27] ) );
  OR2_X1 U76 ( .A1(n93), .A2(n81), .ZN(n80) );
  INV_X1 U78 ( .A(\ab[1][27] ), .ZN(n81) );
  CLKBUF_X3 U80 ( .A(n17), .Z(n82) );
  CLKBUF_X3 U82 ( .A(n63), .Z(n94) );
  CLKBUF_X1 U84 ( .A(n16), .Z(n171) );
  CLKBUF_X3 U85 ( .A(n39), .Z(n106) );
  AND2_X1 U86 ( .A1(B[26]), .A2(A[1]), .ZN(\ab[1][26] ) );
  BUF_X1 U88 ( .A(n15), .Z(n174) );
  AND2_X1 U90 ( .A1(B[29]), .A2(A[2]), .ZN(\ab[2][29] ) );
  AND2_X1 U92 ( .A1(B[27]), .A2(n84), .ZN(\ab[0][27] ) );
  AND2_X1 U94 ( .A1(B[27]), .A2(A[1]), .ZN(\ab[1][27] ) );
  AND2_X1 U96 ( .A1(B[28]), .A2(A[1]), .ZN(\ab[1][28] ) );
  AND2_X1 U98 ( .A1(n63), .A2(ZB), .ZN(\ab[0][31] ) );
  AND2_X1 U100 ( .A1(B[30]), .A2(n84), .ZN(\ab[0][30] ) );
  BUF_X1 U102 ( .A(n12), .Z(n179) );
  CLKBUF_X1 U104 ( .A(n17), .Z(n169) );
  CLKBUF_X1 U106 ( .A(n17), .Z(n167) );
  AND2_X1 U108 ( .A1(B[29]), .A2(A[1]), .ZN(\ab[1][29] ) );
  XOR2_X1 U110 ( .A(\SUMB[31][3] ), .B(\CARRYB[31][2] ), .Z(\A1[32] ) );
  CLKBUF_X1 U112 ( .A(n15), .Z(n175) );
  CLKBUF_X3 U114 ( .A(n15), .Z(n173) );
  CLKBUF_X2 U116 ( .A(QB), .Z(n208) );
  CLKBUF_X2 U118 ( .A(QB), .Z(n209) );
  AND2_X1 U120 ( .A1(B[30]), .A2(A[1]), .ZN(\ab[1][30] ) );
  XNOR2_X1 U122 ( .A(\SUMB[30][2] ), .B(n83), .ZN(\SUMB[31][1] ) );
  XNOR2_X1 U124 ( .A(\CARRYB[30][1] ), .B(\ab[31][1] ), .ZN(n83) );
  XNOR2_X1 U126 ( .A(n85), .B(\ab[0][28] ), .ZN(\SUMB[1][27] ) );
  OR2_X1 U128 ( .A1(n14), .A2(n100), .ZN(n85) );
  BUF_X1 U130 ( .A(n10), .Z(n184) );
  NAND2_X1 U132 ( .A1(\SUMB[30][2] ), .A2(\CARRYB[30][1] ), .ZN(n86) );
  NAND2_X1 U134 ( .A1(\SUMB[30][2] ), .A2(\ab[31][1] ), .ZN(n87) );
  NAND2_X1 U136 ( .A1(\CARRYB[30][1] ), .A2(\ab[31][1] ), .ZN(n88) );
  NAND3_X1 U138 ( .A1(n86), .A2(n87), .A3(n88), .ZN(\CARRYB[31][1] ) );
  INV_X1 U140 ( .A(n184), .ZN(n89) );
  INV_X1 U142 ( .A(n89), .ZN(n91) );
  INV_X1 U144 ( .A(n89), .ZN(n90) );
  CLKBUF_X2 U146 ( .A(n41), .Z(n104) );
  CLKBUF_X3 U148 ( .A(n41), .Z(n105) );
  INV_X1 U150 ( .A(A[1]), .ZN(n92) );
  CLKBUF_X1 U152 ( .A(n35), .Z(n117) );
  BUF_X1 U154 ( .A(n13), .Z(n177) );
  BUF_X1 U156 ( .A(n39), .Z(n107) );
  BUF_X1 U157 ( .A(n38), .Z(n109) );
  BUF_X2 U158 ( .A(n31), .Z(n128) );
  BUF_X2 U160 ( .A(n30), .Z(n131) );
  BUF_X2 U161 ( .A(n26), .Z(n143) );
  BUF_X2 U162 ( .A(n29), .Z(n134) );
  BUF_X2 U164 ( .A(n27), .Z(n140) );
  BUF_X2 U166 ( .A(n25), .Z(n146) );
  BUF_X2 U168 ( .A(n28), .Z(n137) );
  BUF_X2 U170 ( .A(n24), .Z(n149) );
  BUF_X2 U172 ( .A(n24), .Z(n148) );
  BUF_X2 U174 ( .A(n25), .Z(n145) );
  BUF_X1 U176 ( .A(n22), .Z(n155) );
  BUF_X1 U177 ( .A(n33), .Z(n122) );
  BUF_X1 U178 ( .A(n37), .Z(n111) );
  BUF_X1 U180 ( .A(n36), .Z(n113) );
  BUF_X1 U182 ( .A(n35), .Z(n115) );
  BUF_X1 U184 ( .A(n35), .Z(n116) );
  BUF_X1 U186 ( .A(n34), .Z(n118) );
  BUF_X1 U188 ( .A(n34), .Z(n119) );
  BUF_X2 U189 ( .A(n3), .Z(n204) );
  BUF_X2 U190 ( .A(n32), .Z(n125) );
  BUF_X2 U191 ( .A(n9), .Z(n187) );
  BUF_X2 U192 ( .A(n22), .Z(n154) );
  BUF_X2 U193 ( .A(n33), .Z(n121) );
  INV_X1 U194 ( .A(\CARRYB[31][31] ), .ZN(\A1[61] ) );
  NOR2_X1 U195 ( .A1(n179), .A2(n93), .ZN(\ab[0][29] ) );
  NOR2_X1 U196 ( .A1(n13), .A2(n93), .ZN(\ab[0][28] ) );
  NOR2_X1 U197 ( .A1(n171), .A2(n95), .ZN(\ab[0][25] ) );
  NOR2_X1 U198 ( .A1(n168), .A2(n94), .ZN(\ab[0][24] ) );
  NOR2_X1 U199 ( .A1(n18), .A2(n95), .ZN(\ab[0][23] ) );
  NOR2_X1 U200 ( .A1(n162), .A2(n95), .ZN(\ab[0][21] ) );
  NOR2_X1 U201 ( .A1(n19), .A2(n94), .ZN(\ab[0][22] ) );
  NOR2_X1 U202 ( .A1(n159), .A2(n95), .ZN(\ab[0][20] ) );
  NOR2_X1 U203 ( .A1(n153), .A2(n95), .ZN(\ab[0][19] ) );
  NOR2_X1 U204 ( .A1(n150), .A2(n94), .ZN(\ab[0][18] ) );
  NOR2_X1 U205 ( .A1(n147), .A2(n94), .ZN(\ab[0][17] ) );
  NOR2_X1 U206 ( .A1(n144), .A2(n95), .ZN(\ab[0][16] ) );
  NOR2_X1 U207 ( .A1(n141), .A2(n94), .ZN(\ab[0][15] ) );
  NOR2_X1 U208 ( .A1(n135), .A2(n95), .ZN(\ab[0][13] ) );
  NOR2_X1 U209 ( .A1(n138), .A2(n94), .ZN(\ab[0][14] ) );
  NOR2_X1 U210 ( .A1(n132), .A2(n94), .ZN(\ab[0][12] ) );
  NOR2_X1 U211 ( .A1(n129), .A2(n95), .ZN(\ab[0][11] ) );
  NOR2_X1 U212 ( .A1(n126), .A2(n95), .ZN(\ab[0][10] ) );
  NOR2_X1 U213 ( .A1(n205), .A2(n94), .ZN(\ab[0][9] ) );
  NOR2_X1 U214 ( .A1(n202), .A2(n95), .ZN(\ab[0][8] ) );
  NOR2_X1 U215 ( .A1(n199), .A2(n94), .ZN(\ab[0][7] ) );
  NOR2_X1 U216 ( .A1(n196), .A2(n94), .ZN(\ab[0][6] ) );
  NOR2_X1 U217 ( .A1(n193), .A2(n95), .ZN(\ab[0][5] ) );
  NOR2_X1 U218 ( .A1(n190), .A2(n94), .ZN(\ab[0][4] ) );
  NOR2_X1 U219 ( .A1(n183), .A2(n94), .ZN(\ab[0][2] ) );
  NOR2_X1 U220 ( .A1(n188), .A2(n95), .ZN(\ab[0][3] ) );
  NOR2_X1 U221 ( .A1(n156), .A2(n95), .ZN(\ab[0][1] ) );
  NOR2_X1 U222 ( .A1(n140), .A2(n101), .ZN(\ab[1][15] ) );
  NOR2_X1 U223 ( .A1(n137), .A2(n101), .ZN(\ab[1][14] ) );
  NOR2_X1 U224 ( .A1(n134), .A2(n102), .ZN(\ab[1][13] ) );
  NOR2_X1 U225 ( .A1(n131), .A2(n101), .ZN(\ab[1][12] ) );
  NOR2_X1 U226 ( .A1(n128), .A2(n102), .ZN(\ab[1][11] ) );
  NOR2_X1 U227 ( .A1(n125), .A2(n102), .ZN(\ab[1][10] ) );
  NOR2_X1 U228 ( .A1(n122), .A2(n101), .ZN(\ab[1][0] ) );
  NOR2_X1 U229 ( .A1(n171), .A2(n102), .ZN(\ab[1][25] ) );
  NOR2_X1 U230 ( .A1(n168), .A2(n101), .ZN(\ab[1][24] ) );
  NOR2_X1 U231 ( .A1(n166), .A2(n102), .ZN(\ab[1][23] ) );
  NOR2_X1 U232 ( .A1(n19), .A2(n101), .ZN(\ab[1][22] ) );
  NOR2_X1 U233 ( .A1(n161), .A2(n102), .ZN(\ab[1][21] ) );
  NOR2_X1 U234 ( .A1(n158), .A2(n102), .ZN(\ab[1][20] ) );
  NOR2_X1 U235 ( .A1(n152), .A2(n102), .ZN(\ab[1][19] ) );
  NOR2_X1 U236 ( .A1(n149), .A2(n101), .ZN(\ab[1][18] ) );
  NOR2_X1 U237 ( .A1(n146), .A2(n101), .ZN(\ab[1][17] ) );
  NOR2_X1 U238 ( .A1(n143), .A2(n102), .ZN(\ab[1][16] ) );
  NOR2_X1 U239 ( .A1(n201), .A2(n102), .ZN(\ab[1][8] ) );
  NOR2_X1 U240 ( .A1(n204), .A2(n101), .ZN(\ab[1][9] ) );
  NOR2_X1 U241 ( .A1(n198), .A2(n101), .ZN(\ab[1][7] ) );
  NOR2_X1 U242 ( .A1(n195), .A2(n101), .ZN(\ab[1][6] ) );
  NOR2_X1 U243 ( .A1(n192), .A2(n74), .ZN(\ab[1][5] ) );
  NOR2_X1 U244 ( .A1(n8), .A2(n101), .ZN(\ab[1][4] ) );
  NOR2_X1 U245 ( .A1(n182), .A2(n101), .ZN(\ab[1][2] ) );
  NOR2_X1 U246 ( .A1(n187), .A2(n74), .ZN(\ab[1][3] ) );
  NOR2_X1 U247 ( .A1(n155), .A2(n74), .ZN(\ab[1][1] ) );
  NOR2_X1 U248 ( .A1(n103), .A2(n14), .ZN(\ab[2][27] ) );
  NOR2_X1 U249 ( .A1(n13), .A2(n103), .ZN(\ab[2][28] ) );
  AND2_X1 U250 ( .A1(\ab[0][29] ), .A2(\ab[1][28] ), .ZN(\CARRYB[1][28] ) );
  NOR2_X1 U251 ( .A1(n174), .A2(n103), .ZN(\ab[2][26] ) );
  AND2_X1 U252 ( .A1(\ab[1][26] ), .A2(\ab[0][27] ), .ZN(\CARRYB[1][26] ) );
  NOR2_X1 U253 ( .A1(n172), .A2(n105), .ZN(\ab[2][25] ) );
  AND2_X1 U254 ( .A1(\ab[1][25] ), .A2(\ab[0][26] ), .ZN(\CARRYB[1][25] ) );
  NOR2_X1 U255 ( .A1(n82), .A2(n104), .ZN(\ab[2][24] ) );
  AND2_X1 U256 ( .A1(\ab[1][24] ), .A2(\ab[0][25] ), .ZN(\CARRYB[1][24] ) );
  NOR2_X1 U257 ( .A1(n165), .A2(n105), .ZN(\ab[2][23] ) );
  AND2_X1 U258 ( .A1(\ab[1][23] ), .A2(\ab[0][24] ), .ZN(\CARRYB[1][23] ) );
  NOR2_X1 U259 ( .A1(n163), .A2(n104), .ZN(\ab[2][22] ) );
  AND2_X1 U260 ( .A1(\ab[1][22] ), .A2(\ab[0][23] ), .ZN(\CARRYB[1][22] ) );
  NOR2_X1 U261 ( .A1(n160), .A2(n105), .ZN(\ab[2][21] ) );
  AND2_X1 U262 ( .A1(\ab[1][21] ), .A2(\ab[0][22] ), .ZN(\CARRYB[1][21] ) );
  NOR2_X1 U263 ( .A1(n157), .A2(n105), .ZN(\ab[2][20] ) );
  AND2_X1 U264 ( .A1(\ab[1][20] ), .A2(\ab[0][21] ), .ZN(\CARRYB[1][20] ) );
  NOR2_X1 U265 ( .A1(n200), .A2(n105), .ZN(\ab[2][8] ) );
  AND2_X1 U266 ( .A1(\ab[1][8] ), .A2(\ab[0][9] ), .ZN(\CARRYB[1][8] ) );
  NOR2_X1 U267 ( .A1(n191), .A2(n40), .ZN(\ab[30][5] ) );
  NOR2_X1 U268 ( .A1(n186), .A2(n40), .ZN(\ab[30][3] ) );
  NOR2_X1 U269 ( .A1(n181), .A2(n40), .ZN(\ab[30][2] ) );
  NOR2_X1 U270 ( .A1(n194), .A2(n40), .ZN(\ab[30][6] ) );
  NOR2_X1 U271 ( .A1(n186), .A2(n42), .ZN(\ab[29][3] ) );
  NOR2_X1 U272 ( .A1(n194), .A2(n42), .ZN(\ab[29][6] ) );
  NOR2_X1 U273 ( .A1(n136), .A2(n40), .ZN(\ab[30][14] ) );
  NOR2_X1 U274 ( .A1(n189), .A2(n43), .ZN(\ab[28][4] ) );
  NOR2_X1 U275 ( .A1(n194), .A2(n43), .ZN(\ab[28][6] ) );
  NOR2_X1 U276 ( .A1(n197), .A2(n40), .ZN(\ab[30][7] ) );
  NOR2_X1 U277 ( .A1(n133), .A2(n40), .ZN(\ab[30][13] ) );
  NOR2_X1 U278 ( .A1(n139), .A2(n40), .ZN(\ab[30][15] ) );
  NOR2_X1 U279 ( .A1(n154), .A2(n40), .ZN(\ab[30][1] ) );
  NOR2_X1 U280 ( .A1(n181), .A2(n42), .ZN(\ab[29][2] ) );
  NOR2_X1 U281 ( .A1(n197), .A2(n42), .ZN(\ab[29][7] ) );
  NOR2_X1 U282 ( .A1(n203), .A2(n40), .ZN(\ab[30][9] ) );
  NOR2_X1 U283 ( .A1(n186), .A2(n43), .ZN(\ab[28][3] ) );
  NOR2_X1 U284 ( .A1(n191), .A2(n44), .ZN(\ab[27][5] ) );
  NOR2_X1 U285 ( .A1(n194), .A2(n44), .ZN(\ab[27][6] ) );
  NOR2_X1 U286 ( .A1(n197), .A2(n43), .ZN(\ab[28][7] ) );
  NOR2_X1 U287 ( .A1(n130), .A2(n40), .ZN(\ab[30][12] ) );
  NOR2_X1 U288 ( .A1(n124), .A2(n40), .ZN(\ab[30][10] ) );
  NOR2_X1 U289 ( .A1(n136), .A2(n42), .ZN(\ab[29][14] ) );
  NOR2_X1 U290 ( .A1(n139), .A2(n42), .ZN(\ab[29][15] ) );
  NOR2_X1 U291 ( .A1(n189), .A2(n44), .ZN(\ab[27][4] ) );
  NOR2_X1 U292 ( .A1(n127), .A2(n40), .ZN(\ab[30][11] ) );
  NOR2_X1 U293 ( .A1(n197), .A2(n44), .ZN(\ab[27][7] ) );
  NOR2_X1 U294 ( .A1(n195), .A2(n45), .ZN(\ab[26][6] ) );
  NOR2_X1 U295 ( .A1(n133), .A2(n42), .ZN(\ab[29][13] ) );
  NOR2_X1 U296 ( .A1(n192), .A2(n45), .ZN(\ab[26][5] ) );
  NOR2_X1 U297 ( .A1(n124), .A2(n42), .ZN(\ab[29][10] ) );
  NOR2_X1 U298 ( .A1(n200), .A2(n43), .ZN(\ab[28][8] ) );
  NOR2_X1 U299 ( .A1(n181), .A2(n43), .ZN(\ab[28][2] ) );
  NOR2_X1 U300 ( .A1(n127), .A2(n42), .ZN(\ab[29][11] ) );
  NOR2_X1 U301 ( .A1(n200), .A2(n44), .ZN(\ab[27][8] ) );
  NOR2_X1 U302 ( .A1(n139), .A2(n43), .ZN(\ab[28][15] ) );
  NOR2_X1 U303 ( .A1(n189), .A2(n45), .ZN(\ab[26][4] ) );
  NOR2_X1 U304 ( .A1(n136), .A2(n43), .ZN(\ab[28][14] ) );
  NOR2_X1 U305 ( .A1(n195), .A2(n46), .ZN(\ab[25][6] ) );
  NOR2_X1 U306 ( .A1(n201), .A2(n45), .ZN(\ab[26][8] ) );
  NOR2_X1 U307 ( .A1(n124), .A2(n43), .ZN(\ab[28][10] ) );
  NOR2_X1 U308 ( .A1(n198), .A2(n46), .ZN(\ab[25][7] ) );
  NOR2_X1 U309 ( .A1(n142), .A2(n42), .ZN(\ab[29][16] ) );
  NOR2_X1 U310 ( .A1(n127), .A2(n43), .ZN(\ab[28][11] ) );
  NOR2_X1 U311 ( .A1(n142), .A2(n43), .ZN(\ab[28][16] ) );
  NOR2_X1 U312 ( .A1(n192), .A2(n46), .ZN(\ab[25][5] ) );
  NOR2_X1 U313 ( .A1(n203), .A2(n44), .ZN(\ab[27][9] ) );
  NOR2_X1 U314 ( .A1(n133), .A2(n43), .ZN(\ab[28][13] ) );
  NOR2_X1 U315 ( .A1(n130), .A2(n43), .ZN(\ab[28][12] ) );
  NOR2_X1 U316 ( .A1(n201), .A2(n46), .ZN(\ab[25][8] ) );
  NOR2_X1 U317 ( .A1(n139), .A2(n44), .ZN(\ab[27][15] ) );
  NOR2_X1 U318 ( .A1(n124), .A2(n44), .ZN(\ab[27][10] ) );
  NOR2_X1 U319 ( .A1(n204), .A2(n45), .ZN(\ab[26][9] ) );
  NOR2_X1 U320 ( .A1(n198), .A2(n47), .ZN(\ab[24][7] ) );
  NOR2_X1 U321 ( .A1(n142), .A2(n44), .ZN(\ab[27][16] ) );
  NOR2_X1 U322 ( .A1(n195), .A2(n47), .ZN(\ab[24][6] ) );
  NOR2_X1 U323 ( .A1(n142), .A2(n40), .ZN(\ab[30][16] ) );
  NOR2_X1 U324 ( .A1(n136), .A2(n44), .ZN(\ab[27][14] ) );
  NOR2_X1 U325 ( .A1(n201), .A2(n47), .ZN(\ab[24][8] ) );
  NOR2_X1 U326 ( .A1(n181), .A2(n44), .ZN(\ab[27][2] ) );
  NOR2_X1 U327 ( .A1(n189), .A2(n46), .ZN(\ab[25][4] ) );
  NOR2_X1 U328 ( .A1(n204), .A2(n46), .ZN(\ab[25][9] ) );
  NOR2_X1 U329 ( .A1(n130), .A2(n44), .ZN(\ab[27][12] ) );
  NOR2_X1 U330 ( .A1(n133), .A2(n44), .ZN(\ab[27][13] ) );
  NOR2_X1 U331 ( .A1(n125), .A2(n45), .ZN(\ab[26][10] ) );
  NOR2_X1 U332 ( .A1(n204), .A2(n47), .ZN(\ab[24][9] ) );
  NOR2_X1 U333 ( .A1(n201), .A2(n48), .ZN(\ab[23][8] ) );
  NOR2_X1 U334 ( .A1(n143), .A2(n45), .ZN(\ab[26][16] ) );
  NOR2_X1 U335 ( .A1(n140), .A2(n45), .ZN(\ab[26][15] ) );
  NOR2_X1 U336 ( .A1(n125), .A2(n46), .ZN(\ab[25][10] ) );
  NOR2_X1 U337 ( .A1(n131), .A2(n45), .ZN(\ab[26][12] ) );
  NOR2_X1 U338 ( .A1(n195), .A2(n48), .ZN(\ab[23][6] ) );
  NOR2_X1 U339 ( .A1(n137), .A2(n45), .ZN(\ab[26][14] ) );
  NOR2_X1 U340 ( .A1(n145), .A2(n44), .ZN(\ab[27][17] ) );
  NOR2_X1 U341 ( .A1(n134), .A2(n45), .ZN(\ab[26][13] ) );
  NOR2_X1 U342 ( .A1(n204), .A2(n48), .ZN(\ab[23][9] ) );
  NOR2_X1 U343 ( .A1(n125), .A2(n47), .ZN(\ab[24][10] ) );
  NOR2_X1 U344 ( .A1(n145), .A2(n43), .ZN(\ab[28][17] ) );
  NOR2_X1 U345 ( .A1(n128), .A2(n46), .ZN(\ab[25][11] ) );
  NOR2_X1 U346 ( .A1(n146), .A2(n45), .ZN(\ab[26][17] ) );
  NOR2_X1 U347 ( .A1(n189), .A2(n47), .ZN(\ab[24][4] ) );
  NOR2_X1 U348 ( .A1(n201), .A2(n49), .ZN(\ab[22][8] ) );
  NOR2_X1 U349 ( .A1(n131), .A2(n46), .ZN(\ab[25][12] ) );
  NOR2_X1 U350 ( .A1(n204), .A2(n49), .ZN(\ab[22][9] ) );
  NOR2_X1 U351 ( .A1(n125), .A2(n48), .ZN(\ab[23][10] ) );
  NOR2_X1 U352 ( .A1(n143), .A2(n46), .ZN(\ab[25][16] ) );
  NOR2_X1 U353 ( .A1(n182), .A2(n45), .ZN(\ab[26][2] ) );
  NOR2_X1 U354 ( .A1(n140), .A2(n46), .ZN(\ab[25][15] ) );
  NOR2_X1 U355 ( .A1(n134), .A2(n46), .ZN(\ab[25][13] ) );
  NOR2_X1 U356 ( .A1(n128), .A2(n47), .ZN(\ab[24][11] ) );
  NOR2_X1 U357 ( .A1(n137), .A2(n46), .ZN(\ab[25][14] ) );
  NOR2_X1 U358 ( .A1(n146), .A2(n46), .ZN(\ab[25][17] ) );
  NOR2_X1 U359 ( .A1(n195), .A2(n49), .ZN(\ab[22][6] ) );
  NOR2_X1 U360 ( .A1(n125), .A2(n49), .ZN(\ab[22][10] ) );
  NOR2_X1 U361 ( .A1(n145), .A2(n42), .ZN(\ab[29][17] ) );
  NOR2_X1 U362 ( .A1(n131), .A2(n47), .ZN(\ab[24][12] ) );
  NOR2_X1 U363 ( .A1(n201), .A2(n50), .ZN(\ab[21][8] ) );
  NOR2_X1 U364 ( .A1(n143), .A2(n47), .ZN(\ab[24][16] ) );
  NOR2_X1 U365 ( .A1(n125), .A2(n50), .ZN(\ab[21][10] ) );
  NOR2_X1 U366 ( .A1(n140), .A2(n47), .ZN(\ab[24][15] ) );
  NOR2_X1 U367 ( .A1(n137), .A2(n47), .ZN(\ab[24][14] ) );
  NOR2_X1 U368 ( .A1(n146), .A2(n47), .ZN(\ab[24][17] ) );
  NOR2_X1 U369 ( .A1(n189), .A2(n48), .ZN(\ab[23][4] ) );
  NOR2_X1 U370 ( .A1(n149), .A2(n45), .ZN(\ab[26][18] ) );
  NOR2_X1 U371 ( .A1(n131), .A2(n48), .ZN(\ab[23][12] ) );
  NOR2_X1 U372 ( .A1(n149), .A2(n46), .ZN(\ab[25][18] ) );
  NOR2_X1 U373 ( .A1(n148), .A2(n44), .ZN(\ab[27][18] ) );
  NOR2_X1 U374 ( .A1(n201), .A2(n51), .ZN(\ab[20][8] ) );
  NOR2_X1 U375 ( .A1(n195), .A2(n50), .ZN(\ab[21][6] ) );
  NOR2_X1 U376 ( .A1(n128), .A2(n50), .ZN(\ab[21][11] ) );
  NOR2_X1 U377 ( .A1(n134), .A2(n48), .ZN(\ab[23][13] ) );
  NOR2_X1 U378 ( .A1(n125), .A2(n51), .ZN(\ab[20][10] ) );
  NOR2_X1 U379 ( .A1(n148), .A2(n43), .ZN(\ab[28][18] ) );
  NOR2_X1 U380 ( .A1(n149), .A2(n47), .ZN(\ab[24][18] ) );
  NOR2_X1 U381 ( .A1(n131), .A2(n49), .ZN(\ab[22][12] ) );
  NOR2_X1 U382 ( .A1(n182), .A2(n46), .ZN(\ab[25][2] ) );
  NOR2_X1 U383 ( .A1(n137), .A2(n48), .ZN(\ab[23][14] ) );
  NOR2_X1 U384 ( .A1(n143), .A2(n48), .ZN(\ab[23][16] ) );
  NOR2_X1 U385 ( .A1(n146), .A2(n48), .ZN(\ab[23][17] ) );
  NOR2_X1 U386 ( .A1(n128), .A2(n51), .ZN(\ab[20][11] ) );
  NOR2_X1 U387 ( .A1(n131), .A2(n50), .ZN(\ab[21][12] ) );
  NOR2_X1 U388 ( .A1(n134), .A2(n49), .ZN(\ab[22][13] ) );
  NOR2_X1 U389 ( .A1(n151), .A2(n44), .ZN(\ab[27][19] ) );
  NOR2_X1 U390 ( .A1(n125), .A2(n53), .ZN(\ab[19][10] ) );
  NOR2_X1 U391 ( .A1(n149), .A2(n48), .ZN(\ab[23][18] ) );
  NOR2_X1 U392 ( .A1(n201), .A2(n53), .ZN(\ab[19][8] ) );
  NOR2_X1 U393 ( .A1(n137), .A2(n49), .ZN(\ab[22][14] ) );
  NOR2_X1 U394 ( .A1(n189), .A2(n49), .ZN(\ab[22][4] ) );
  NOR2_X1 U395 ( .A1(n131), .A2(n51), .ZN(\ab[20][12] ) );
  NOR2_X1 U396 ( .A1(n158), .A2(n45), .ZN(\ab[26][20] ) );
  NOR2_X1 U397 ( .A1(n143), .A2(n49), .ZN(\ab[22][16] ) );
  NOR2_X1 U398 ( .A1(n195), .A2(n51), .ZN(\ab[20][6] ) );
  NOR2_X1 U399 ( .A1(n146), .A2(n49), .ZN(\ab[22][17] ) );
  NOR2_X1 U400 ( .A1(n152), .A2(n45), .ZN(\ab[26][19] ) );
  NOR2_X1 U401 ( .A1(n152), .A2(n46), .ZN(\ab[25][19] ) );
  NOR2_X1 U402 ( .A1(n152), .A2(n47), .ZN(\ab[24][19] ) );
  NOR2_X1 U403 ( .A1(n125), .A2(n54), .ZN(\ab[18][10] ) );
  NOR2_X1 U404 ( .A1(n149), .A2(n49), .ZN(\ab[22][18] ) );
  NOR2_X1 U405 ( .A1(n131), .A2(n53), .ZN(\ab[19][12] ) );
  NOR2_X1 U406 ( .A1(n137), .A2(n50), .ZN(\ab[21][14] ) );
  NOR2_X1 U407 ( .A1(n152), .A2(n48), .ZN(\ab[23][19] ) );
  NOR2_X1 U408 ( .A1(n161), .A2(n46), .ZN(\ab[25][21] ) );
  NOR2_X1 U409 ( .A1(n140), .A2(n50), .ZN(\ab[21][15] ) );
  NOR2_X1 U410 ( .A1(n182), .A2(n47), .ZN(\ab[24][2] ) );
  NOR2_X1 U411 ( .A1(n201), .A2(n54), .ZN(\ab[18][8] ) );
  NOR2_X1 U412 ( .A1(n143), .A2(n50), .ZN(\ab[21][16] ) );
  NOR2_X1 U413 ( .A1(n131), .A2(n54), .ZN(\ab[18][12] ) );
  NOR2_X1 U414 ( .A1(n152), .A2(n49), .ZN(\ab[22][19] ) );
  NOR2_X1 U415 ( .A1(n134), .A2(n53), .ZN(\ab[19][13] ) );
  NOR2_X1 U416 ( .A1(n137), .A2(n51), .ZN(\ab[20][14] ) );
  NOR2_X1 U417 ( .A1(n149), .A2(n50), .ZN(\ab[21][18] ) );
  NOR2_X1 U418 ( .A1(n158), .A2(n46), .ZN(\ab[25][20] ) );
  NOR2_X1 U419 ( .A1(n125), .A2(n55), .ZN(\ab[17][10] ) );
  NOR2_X1 U420 ( .A1(n195), .A2(n53), .ZN(\ab[19][6] ) );
  NOR2_X1 U421 ( .A1(n189), .A2(n50), .ZN(\ab[21][4] ) );
  NOR2_X1 U422 ( .A1(n140), .A2(n51), .ZN(\ab[20][15] ) );
  NOR2_X1 U423 ( .A1(n131), .A2(n55), .ZN(\ab[17][12] ) );
  NOR2_X1 U424 ( .A1(n134), .A2(n54), .ZN(\ab[18][13] ) );
  NOR2_X1 U425 ( .A1(n163), .A2(n47), .ZN(\ab[24][22] ) );
  NOR2_X1 U426 ( .A1(n152), .A2(n50), .ZN(\ab[21][19] ) );
  NOR2_X1 U427 ( .A1(n158), .A2(n47), .ZN(\ab[24][20] ) );
  NOR2_X1 U428 ( .A1(n137), .A2(n53), .ZN(\ab[19][14] ) );
  NOR2_X1 U429 ( .A1(n143), .A2(n51), .ZN(\ab[20][16] ) );
  NOR2_X1 U430 ( .A1(n158), .A2(n48), .ZN(\ab[23][20] ) );
  NOR2_X1 U431 ( .A1(n149), .A2(n51), .ZN(\ab[20][18] ) );
  NOR2_X1 U432 ( .A1(n158), .A2(n49), .ZN(\ab[22][20] ) );
  NOR2_X1 U433 ( .A1(n201), .A2(n55), .ZN(\ab[17][8] ) );
  NOR2_X1 U434 ( .A1(n161), .A2(n47), .ZN(\ab[24][21] ) );
  NOR2_X1 U435 ( .A1(n125), .A2(n56), .ZN(\ab[16][10] ) );
  NOR2_X1 U436 ( .A1(n137), .A2(n54), .ZN(\ab[18][14] ) );
  NOR2_X1 U437 ( .A1(n131), .A2(n56), .ZN(\ab[16][12] ) );
  NOR2_X1 U438 ( .A1(n152), .A2(n51), .ZN(\ab[20][19] ) );
  NOR2_X1 U439 ( .A1(n182), .A2(n48), .ZN(\ab[23][2] ) );
  NOR2_X1 U440 ( .A1(n143), .A2(n53), .ZN(\ab[19][16] ) );
  NOR2_X1 U441 ( .A1(n158), .A2(n50), .ZN(\ab[21][20] ) );
  NOR2_X1 U442 ( .A1(n192), .A2(n53), .ZN(\ab[19][5] ) );
  NOR2_X1 U443 ( .A1(n146), .A2(n53), .ZN(\ab[19][17] ) );
  NOR2_X1 U444 ( .A1(n137), .A2(n55), .ZN(\ab[17][14] ) );
  NOR2_X1 U445 ( .A1(n73), .A2(n48), .ZN(\ab[23][23] ) );
  NOR2_X1 U446 ( .A1(n149), .A2(n53), .ZN(\ab[19][18] ) );
  NOR2_X1 U447 ( .A1(n198), .A2(n55), .ZN(\ab[17][7] ) );
  NOR2_X1 U448 ( .A1(n187), .A2(n50), .ZN(\ab[21][3] ) );
  NOR2_X1 U449 ( .A1(n161), .A2(n48), .ZN(\ab[23][21] ) );
  NOR2_X1 U450 ( .A1(n158), .A2(n51), .ZN(\ab[20][20] ) );
  NOR2_X1 U451 ( .A1(n164), .A2(n48), .ZN(\ab[23][22] ) );
  NOR2_X1 U452 ( .A1(n132), .A2(n57), .ZN(\ab[15][12] ) );
  NOR2_X1 U453 ( .A1(n137), .A2(n56), .ZN(\ab[16][14] ) );
  NOR2_X1 U454 ( .A1(n152), .A2(n53), .ZN(\ab[19][19] ) );
  NOR2_X1 U455 ( .A1(n143), .A2(n54), .ZN(\ab[18][16] ) );
  NOR2_X1 U456 ( .A1(n140), .A2(n55), .ZN(\ab[17][15] ) );
  NOR2_X1 U457 ( .A1(n176), .A2(n109), .ZN(\ab[4][27] ) );
  NOR2_X1 U458 ( .A1(n170), .A2(n114), .ZN(\ab[6][25] ) );
  NOR2_X1 U459 ( .A1(n165), .A2(n119), .ZN(\ab[8][23] ) );
  NOR2_X1 U460 ( .A1(n162), .A2(n96), .ZN(\ab[10][21] ) );
  NOR2_X1 U461 ( .A1(n153), .A2(n98), .ZN(\ab[12][19] ) );
  NOR2_X1 U462 ( .A1(n147), .A2(n58), .ZN(\ab[14][17] ) );
  NOR2_X1 U463 ( .A1(n140), .A2(n56), .ZN(\ab[16][15] ) );
  NOR2_X1 U464 ( .A1(n177), .A2(n106), .ZN(\ab[3][28] ) );
  NOR2_X1 U465 ( .A1(n175), .A2(n112), .ZN(\ab[5][26] ) );
  NOR2_X1 U466 ( .A1(n167), .A2(n116), .ZN(\ab[7][24] ) );
  NOR2_X1 U467 ( .A1(n207), .A2(n164), .ZN(\ab[9][22] ) );
  NOR2_X1 U468 ( .A1(n159), .A2(n97), .ZN(\ab[11][20] ) );
  NOR2_X1 U469 ( .A1(n150), .A2(n59), .ZN(\ab[13][18] ) );
  NOR2_X1 U470 ( .A1(n144), .A2(n57), .ZN(\ab[15][16] ) );
  NOR2_X1 U471 ( .A1(n176), .A2(n111), .ZN(\ab[5][27] ) );
  NOR2_X1 U472 ( .A1(n170), .A2(n116), .ZN(\ab[7][25] ) );
  NOR2_X1 U473 ( .A1(n207), .A2(n165), .ZN(\ab[9][23] ) );
  NOR2_X1 U474 ( .A1(n162), .A2(n97), .ZN(\ab[11][21] ) );
  NOR2_X1 U475 ( .A1(n153), .A2(n59), .ZN(\ab[13][19] ) );
  NOR2_X1 U476 ( .A1(n147), .A2(n57), .ZN(\ab[15][17] ) );
  NOR2_X1 U477 ( .A1(n170), .A2(n110), .ZN(\ab[4][25] ) );
  NOR2_X1 U478 ( .A1(n170), .A2(n112), .ZN(\ab[5][25] ) );
  NOR2_X1 U479 ( .A1(n165), .A2(n114), .ZN(\ab[6][23] ) );
  NOR2_X1 U480 ( .A1(n165), .A2(n116), .ZN(\ab[7][23] ) );
  NOR2_X1 U481 ( .A1(n176), .A2(n106), .ZN(\ab[3][27] ) );
  NOR2_X1 U482 ( .A1(n175), .A2(n114), .ZN(\ab[6][26] ) );
  NOR2_X1 U483 ( .A1(n169), .A2(n119), .ZN(\ab[8][24] ) );
  NOR2_X1 U484 ( .A1(n163), .A2(n62), .ZN(\ab[10][22] ) );
  NOR2_X1 U485 ( .A1(n159), .A2(n98), .ZN(\ab[12][20] ) );
  NOR2_X1 U486 ( .A1(n150), .A2(n58), .ZN(\ab[14][18] ) );
  NOR2_X1 U487 ( .A1(n143), .A2(n56), .ZN(\ab[16][16] ) );
  NOR2_X1 U488 ( .A1(n177), .A2(n109), .ZN(\ab[4][28] ) );
  NOR2_X1 U489 ( .A1(n176), .A2(n113), .ZN(\ab[6][27] ) );
  NOR2_X1 U490 ( .A1(n73), .A2(n62), .ZN(\ab[10][23] ) );
  NOR2_X1 U491 ( .A1(n176), .A2(n115), .ZN(\ab[7][27] ) );
  NOR2_X1 U492 ( .A1(n173), .A2(n110), .ZN(\ab[4][26] ) );
  NOR2_X1 U493 ( .A1(n82), .A2(n114), .ZN(\ab[6][24] ) );
  NOR2_X1 U494 ( .A1(n163), .A2(n119), .ZN(\ab[8][22] ) );
  NOR2_X1 U495 ( .A1(n159), .A2(n96), .ZN(\ab[10][20] ) );
  NOR2_X1 U496 ( .A1(n150), .A2(n98), .ZN(\ab[12][18] ) );
  NOR2_X1 U497 ( .A1(n144), .A2(n58), .ZN(\ab[14][16] ) );
  NOR2_X1 U498 ( .A1(n207), .A2(n82), .ZN(\ab[9][24] ) );
  NOR2_X1 U499 ( .A1(n163), .A2(n97), .ZN(\ab[11][22] ) );
  NOR2_X1 U500 ( .A1(n164), .A2(n98), .ZN(\ab[12][22] ) );
  NOR2_X1 U501 ( .A1(n159), .A2(n59), .ZN(\ab[13][20] ) );
  NOR2_X1 U502 ( .A1(n159), .A2(n58), .ZN(\ab[14][20] ) );
  NOR2_X1 U503 ( .A1(n150), .A2(n57), .ZN(\ab[15][18] ) );
  NOR2_X1 U504 ( .A1(n149), .A2(n56), .ZN(\ab[16][18] ) );
  NOR2_X1 U505 ( .A1(n143), .A2(n55), .ZN(\ab[17][16] ) );
  NOR2_X1 U506 ( .A1(n173), .A2(n116), .ZN(\ab[7][26] ) );
  NOR2_X1 U507 ( .A1(n82), .A2(n62), .ZN(\ab[10][24] ) );
  NOR2_X1 U508 ( .A1(n178), .A2(n111), .ZN(\ab[5][28] ) );
  NOR2_X1 U509 ( .A1(n175), .A2(n119), .ZN(\ab[8][26] ) );
  NOR2_X1 U510 ( .A1(n177), .A2(n113), .ZN(\ab[6][28] ) );
  NOR2_X1 U511 ( .A1(n126), .A2(n57), .ZN(\ab[15][10] ) );
  NOR2_X1 U512 ( .A1(n173), .A2(n107), .ZN(\ab[3][26] ) );
  NOR2_X1 U513 ( .A1(n82), .A2(n112), .ZN(\ab[5][24] ) );
  NOR2_X1 U514 ( .A1(n163), .A2(n116), .ZN(\ab[7][22] ) );
  NOR2_X1 U515 ( .A1(n207), .A2(n157), .ZN(\ab[9][20] ) );
  NOR2_X1 U516 ( .A1(n150), .A2(n97), .ZN(\ab[11][18] ) );
  NOR2_X1 U517 ( .A1(n144), .A2(n59), .ZN(\ab[13][16] ) );
  NOR2_X1 U518 ( .A1(n138), .A2(n57), .ZN(\ab[15][14] ) );
  NOR2_X1 U519 ( .A1(n159), .A2(n57), .ZN(\ab[15][20] ) );
  NOR2_X1 U520 ( .A1(n149), .A2(n55), .ZN(\ab[17][18] ) );
  NOR2_X1 U521 ( .A1(n163), .A2(n59), .ZN(\ab[13][22] ) );
  NOR2_X1 U522 ( .A1(n82), .A2(n97), .ZN(\ab[11][24] ) );
  NOR2_X1 U523 ( .A1(n207), .A2(n173), .ZN(\ab[9][26] ) );
  NOR2_X1 U524 ( .A1(n178), .A2(n115), .ZN(\ab[7][28] ) );
  NOR2_X1 U525 ( .A1(n161), .A2(n49), .ZN(\ab[22][21] ) );
  NOR2_X1 U526 ( .A1(n73), .A2(n98), .ZN(\ab[12][23] ) );
  NOR2_X1 U527 ( .A1(n162), .A2(n99), .ZN(\ab[14][21] ) );
  NOR2_X1 U528 ( .A1(n152), .A2(n56), .ZN(\ab[16][19] ) );
  NOR2_X1 U529 ( .A1(n146), .A2(n54), .ZN(\ab[18][17] ) );
  NOR2_X1 U530 ( .A1(n172), .A2(n62), .ZN(\ab[10][25] ) );
  NOR2_X1 U531 ( .A1(n176), .A2(n118), .ZN(\ab[8][27] ) );
  NOR2_X1 U532 ( .A1(n169), .A2(n110), .ZN(\ab[4][24] ) );
  NOR2_X1 U533 ( .A1(n164), .A2(n114), .ZN(\ab[6][22] ) );
  NOR2_X1 U534 ( .A1(n157), .A2(n119), .ZN(\ab[8][20] ) );
  NOR2_X1 U535 ( .A1(n150), .A2(n96), .ZN(\ab[10][18] ) );
  NOR2_X1 U536 ( .A1(n144), .A2(n98), .ZN(\ab[12][16] ) );
  NOR2_X1 U537 ( .A1(n138), .A2(n99), .ZN(\ab[14][14] ) );
  NOR2_X1 U538 ( .A1(n152), .A2(n55), .ZN(\ab[17][19] ) );
  NOR2_X1 U539 ( .A1(n162), .A2(n57), .ZN(\ab[15][21] ) );
  NOR2_X1 U540 ( .A1(n73), .A2(n59), .ZN(\ab[13][23] ) );
  NOR2_X1 U541 ( .A1(n170), .A2(n97), .ZN(\ab[11][25] ) );
  NOR2_X1 U542 ( .A1(n206), .A2(n176), .ZN(\ab[9][27] ) );
  NOR2_X1 U543 ( .A1(n149), .A2(n54), .ZN(\ab[18][18] ) );
  NOR2_X1 U544 ( .A1(n158), .A2(n56), .ZN(\ab[16][20] ) );
  NOR2_X1 U545 ( .A1(n163), .A2(n58), .ZN(\ab[14][22] ) );
  NOR2_X1 U546 ( .A1(n82), .A2(n98), .ZN(\ab[12][24] ) );
  NOR2_X1 U547 ( .A1(n175), .A2(n62), .ZN(\ab[10][26] ) );
  NOR2_X1 U548 ( .A1(n178), .A2(n118), .ZN(\ab[8][28] ) );
  NOR2_X1 U549 ( .A1(n165), .A2(n110), .ZN(\ab[4][23] ) );
  NOR2_X1 U550 ( .A1(n167), .A2(n107), .ZN(\ab[3][24] ) );
  NOR2_X1 U551 ( .A1(n163), .A2(n112), .ZN(\ab[5][22] ) );
  NOR2_X1 U552 ( .A1(n157), .A2(n116), .ZN(\ab[7][20] ) );
  NOR2_X1 U553 ( .A1(n207), .A2(n148), .ZN(\ab[9][18] ) );
  NOR2_X1 U554 ( .A1(n144), .A2(n97), .ZN(\ab[11][16] ) );
  NOR2_X1 U555 ( .A1(n138), .A2(n59), .ZN(\ab[13][14] ) );
  NOR2_X1 U556 ( .A1(n161), .A2(n56), .ZN(\ab[16][21] ) );
  NOR2_X1 U557 ( .A1(n73), .A2(n58), .ZN(\ab[14][23] ) );
  NOR2_X1 U558 ( .A1(n161), .A2(n55), .ZN(\ab[17][21] ) );
  NOR2_X1 U559 ( .A1(n170), .A2(n98), .ZN(\ab[12][25] ) );
  NOR2_X1 U560 ( .A1(n73), .A2(n57), .ZN(\ab[15][23] ) );
  NOR2_X1 U561 ( .A1(n176), .A2(n62), .ZN(\ab[10][27] ) );
  NOR2_X1 U562 ( .A1(n170), .A2(n59), .ZN(\ab[13][25] ) );
  NOR2_X1 U563 ( .A1(n176), .A2(n61), .ZN(\ab[11][27] ) );
  NOR2_X1 U564 ( .A1(n158), .A2(n55), .ZN(\ab[17][20] ) );
  NOR2_X1 U565 ( .A1(n163), .A2(n57), .ZN(\ab[15][22] ) );
  NOR2_X1 U566 ( .A1(n158), .A2(n54), .ZN(\ab[18][20] ) );
  NOR2_X1 U567 ( .A1(n167), .A2(n59), .ZN(\ab[13][24] ) );
  NOR2_X1 U568 ( .A1(n163), .A2(n56), .ZN(\ab[16][22] ) );
  NOR2_X1 U569 ( .A1(n173), .A2(n97), .ZN(\ab[11][26] ) );
  NOR2_X1 U570 ( .A1(n169), .A2(n58), .ZN(\ab[14][24] ) );
  NOR2_X1 U571 ( .A1(n206), .A2(n177), .ZN(\ab[9][28] ) );
  NOR2_X1 U572 ( .A1(n173), .A2(n98), .ZN(\ab[12][26] ) );
  NOR2_X1 U573 ( .A1(n178), .A2(n62), .ZN(\ab[10][28] ) );
  NOR2_X1 U574 ( .A1(n164), .A2(n110), .ZN(\ab[4][22] ) );
  NOR2_X1 U575 ( .A1(n157), .A2(n114), .ZN(\ab[6][20] ) );
  NOR2_X1 U576 ( .A1(n148), .A2(n119), .ZN(\ab[8][18] ) );
  NOR2_X1 U577 ( .A1(n144), .A2(n96), .ZN(\ab[10][16] ) );
  NOR2_X1 U578 ( .A1(n138), .A2(n98), .ZN(\ab[12][14] ) );
  NOR2_X1 U579 ( .A1(n132), .A2(n99), .ZN(\ab[14][12] ) );
  NOR2_X1 U580 ( .A1(n158), .A2(n53), .ZN(\ab[19][20] ) );
  NOR2_X1 U581 ( .A1(n164), .A2(n55), .ZN(\ab[17][22] ) );
  NOR2_X1 U582 ( .A1(n82), .A2(n57), .ZN(\ab[15][24] ) );
  NOR2_X1 U583 ( .A1(n175), .A2(n59), .ZN(\ab[13][26] ) );
  NOR2_X1 U584 ( .A1(n178), .A2(n61), .ZN(\ab[11][28] ) );
  NOR2_X1 U585 ( .A1(n161), .A2(n54), .ZN(\ab[18][21] ) );
  NOR2_X1 U586 ( .A1(n73), .A2(n56), .ZN(\ab[16][23] ) );
  NOR2_X1 U587 ( .A1(n172), .A2(n58), .ZN(\ab[14][25] ) );
  NOR2_X1 U588 ( .A1(n176), .A2(n60), .ZN(\ab[12][27] ) );
  NOR2_X1 U589 ( .A1(n164), .A2(n107), .ZN(\ab[3][22] ) );
  NOR2_X1 U590 ( .A1(n157), .A2(n112), .ZN(\ab[5][20] ) );
  NOR2_X1 U591 ( .A1(n148), .A2(n116), .ZN(\ab[7][18] ) );
  NOR2_X1 U592 ( .A1(n207), .A2(n142), .ZN(\ab[9][16] ) );
  NOR2_X1 U593 ( .A1(n138), .A2(n97), .ZN(\ab[11][14] ) );
  NOR2_X1 U594 ( .A1(n132), .A2(n59), .ZN(\ab[13][12] ) );
  NOR2_X1 U595 ( .A1(n161), .A2(n50), .ZN(\ab[21][21] ) );
  NOR2_X1 U596 ( .A1(n160), .A2(n107), .ZN(\ab[3][21] ) );
  NOR2_X1 U597 ( .A1(n151), .A2(n112), .ZN(\ab[5][19] ) );
  NOR2_X1 U598 ( .A1(n145), .A2(n116), .ZN(\ab[7][17] ) );
  NOR2_X1 U599 ( .A1(n207), .A2(n139), .ZN(\ab[9][15] ) );
  NOR2_X1 U600 ( .A1(n135), .A2(n97), .ZN(\ab[11][13] ) );
  NOR2_X1 U601 ( .A1(n129), .A2(n59), .ZN(\ab[13][11] ) );
  NOR2_X1 U602 ( .A1(n205), .A2(n57), .ZN(\ab[15][9] ) );
  NOR2_X1 U603 ( .A1(n155), .A2(n48), .ZN(\ab[23][1] ) );
  NOR2_X1 U604 ( .A1(n148), .A2(n112), .ZN(\ab[5][18] ) );
  NOR2_X1 U605 ( .A1(n157), .A2(n107), .ZN(\ab[3][20] ) );
  NOR2_X1 U606 ( .A1(n142), .A2(n116), .ZN(\ab[7][16] ) );
  NOR2_X1 U607 ( .A1(n207), .A2(n136), .ZN(\ab[9][14] ) );
  NOR2_X1 U608 ( .A1(n132), .A2(n97), .ZN(\ab[11][12] ) );
  NOR2_X1 U609 ( .A1(n126), .A2(n59), .ZN(\ab[13][10] ) );
  NOR2_X1 U610 ( .A1(n202), .A2(n57), .ZN(\ab[15][8] ) );
  NOR2_X1 U611 ( .A1(n195), .A2(n55), .ZN(\ab[17][6] ) );
  NOR2_X1 U612 ( .A1(n189), .A2(n53), .ZN(\ab[19][4] ) );
  NOR2_X1 U613 ( .A1(n182), .A2(n50), .ZN(\ab[21][2] ) );
  NOR2_X1 U614 ( .A1(n151), .A2(n107), .ZN(\ab[3][19] ) );
  NOR2_X1 U615 ( .A1(n145), .A2(n112), .ZN(\ab[5][17] ) );
  NOR2_X1 U616 ( .A1(n139), .A2(n117), .ZN(\ab[7][15] ) );
  NOR2_X1 U617 ( .A1(n207), .A2(n133), .ZN(\ab[9][13] ) );
  NOR2_X1 U618 ( .A1(n129), .A2(n97), .ZN(\ab[11][11] ) );
  NOR2_X1 U619 ( .A1(n205), .A2(n59), .ZN(\ab[13][9] ) );
  NOR2_X1 U620 ( .A1(n199), .A2(n57), .ZN(\ab[15][7] ) );
  NOR2_X1 U621 ( .A1(n192), .A2(n55), .ZN(\ab[17][5] ) );
  NOR2_X1 U622 ( .A1(n187), .A2(n53), .ZN(\ab[19][3] ) );
  NOR2_X1 U623 ( .A1(n155), .A2(n50), .ZN(\ab[21][1] ) );
  NOR2_X1 U624 ( .A1(n148), .A2(n107), .ZN(\ab[3][18] ) );
  NOR2_X1 U625 ( .A1(n142), .A2(n112), .ZN(\ab[5][16] ) );
  NOR2_X1 U626 ( .A1(n136), .A2(n117), .ZN(\ab[7][14] ) );
  NOR2_X1 U627 ( .A1(n207), .A2(n130), .ZN(\ab[9][12] ) );
  NOR2_X1 U628 ( .A1(n126), .A2(n61), .ZN(\ab[11][10] ) );
  NOR2_X1 U629 ( .A1(n202), .A2(n59), .ZN(\ab[13][8] ) );
  NOR2_X1 U630 ( .A1(n196), .A2(n57), .ZN(\ab[15][6] ) );
  NOR2_X1 U631 ( .A1(n189), .A2(n55), .ZN(\ab[17][4] ) );
  NOR2_X1 U632 ( .A1(n182), .A2(n53), .ZN(\ab[19][2] ) );
  NOR2_X1 U633 ( .A1(n163), .A2(n54), .ZN(\ab[18][22] ) );
  NOR2_X1 U634 ( .A1(n82), .A2(n56), .ZN(\ab[16][24] ) );
  NOR2_X1 U635 ( .A1(n173), .A2(n58), .ZN(\ab[14][26] ) );
  NOR2_X1 U636 ( .A1(n177), .A2(n60), .ZN(\ab[12][28] ) );
  NOR2_X1 U637 ( .A1(n161), .A2(n53), .ZN(\ab[19][21] ) );
  NOR2_X1 U638 ( .A1(n73), .A2(n55), .ZN(\ab[17][23] ) );
  NOR2_X1 U639 ( .A1(n170), .A2(n57), .ZN(\ab[15][25] ) );
  NOR2_X1 U640 ( .A1(n176), .A2(n59), .ZN(\ab[13][27] ) );
  NOR2_X1 U641 ( .A1(n145), .A2(n107), .ZN(\ab[3][17] ) );
  NOR2_X1 U642 ( .A1(n139), .A2(n112), .ZN(\ab[5][15] ) );
  NOR2_X1 U643 ( .A1(n133), .A2(n117), .ZN(\ab[7][13] ) );
  NOR2_X1 U644 ( .A1(n207), .A2(n127), .ZN(\ab[9][11] ) );
  NOR2_X1 U645 ( .A1(n205), .A2(n61), .ZN(\ab[11][9] ) );
  NOR2_X1 U646 ( .A1(n199), .A2(n59), .ZN(\ab[13][7] ) );
  NOR2_X1 U647 ( .A1(n193), .A2(n57), .ZN(\ab[15][5] ) );
  NOR2_X1 U648 ( .A1(n187), .A2(n55), .ZN(\ab[17][3] ) );
  NOR2_X1 U649 ( .A1(n155), .A2(n53), .ZN(\ab[19][1] ) );
  NOR2_X1 U650 ( .A1(n142), .A2(n107), .ZN(\ab[3][16] ) );
  NOR2_X1 U651 ( .A1(n136), .A2(n112), .ZN(\ab[5][14] ) );
  NOR2_X1 U652 ( .A1(n130), .A2(n117), .ZN(\ab[7][12] ) );
  NOR2_X1 U653 ( .A1(n207), .A2(n124), .ZN(\ab[9][10] ) );
  NOR2_X1 U654 ( .A1(n202), .A2(n61), .ZN(\ab[11][8] ) );
  NOR2_X1 U655 ( .A1(n196), .A2(n59), .ZN(\ab[13][6] ) );
  NOR2_X1 U656 ( .A1(n190), .A2(n57), .ZN(\ab[15][4] ) );
  NOR2_X1 U657 ( .A1(n182), .A2(n55), .ZN(\ab[17][2] ) );
  NOR2_X1 U658 ( .A1(n163), .A2(n53), .ZN(\ab[19][22] ) );
  NOR2_X1 U659 ( .A1(n167), .A2(n55), .ZN(\ab[17][24] ) );
  NOR2_X1 U660 ( .A1(n173), .A2(n57), .ZN(\ab[15][26] ) );
  NOR2_X1 U661 ( .A1(n178), .A2(n59), .ZN(\ab[13][28] ) );
  NOR2_X1 U662 ( .A1(n161), .A2(n51), .ZN(\ab[20][21] ) );
  NOR2_X1 U663 ( .A1(n73), .A2(n54), .ZN(\ab[18][23] ) );
  NOR2_X1 U664 ( .A1(n170), .A2(n56), .ZN(\ab[16][25] ) );
  NOR2_X1 U665 ( .A1(n73), .A2(n53), .ZN(\ab[19][23] ) );
  NOR2_X1 U666 ( .A1(n176), .A2(n58), .ZN(\ab[14][27] ) );
  NOR2_X1 U667 ( .A1(n170), .A2(n55), .ZN(\ab[17][25] ) );
  NOR2_X1 U668 ( .A1(n176), .A2(n57), .ZN(\ab[15][27] ) );
  NOR2_X1 U669 ( .A1(n139), .A2(n108), .ZN(\ab[3][15] ) );
  NOR2_X1 U670 ( .A1(n133), .A2(n112), .ZN(\ab[5][13] ) );
  NOR2_X1 U671 ( .A1(n127), .A2(n117), .ZN(\ab[7][11] ) );
  NOR2_X1 U672 ( .A1(n206), .A2(n203), .ZN(\ab[9][9] ) );
  NOR2_X1 U673 ( .A1(n199), .A2(n61), .ZN(\ab[11][7] ) );
  NOR2_X1 U674 ( .A1(n193), .A2(n59), .ZN(\ab[13][5] ) );
  NOR2_X1 U675 ( .A1(n188), .A2(n57), .ZN(\ab[15][3] ) );
  NOR2_X1 U676 ( .A1(n155), .A2(n55), .ZN(\ab[17][1] ) );
  NOR2_X1 U677 ( .A1(n164), .A2(n51), .ZN(\ab[20][22] ) );
  NOR2_X1 U678 ( .A1(n169), .A2(n54), .ZN(\ab[18][24] ) );
  NOR2_X1 U679 ( .A1(n173), .A2(n56), .ZN(\ab[16][26] ) );
  NOR2_X1 U680 ( .A1(n178), .A2(n99), .ZN(\ab[14][28] ) );
  NOR2_X1 U681 ( .A1(n163), .A2(n50), .ZN(\ab[21][22] ) );
  NOR2_X1 U682 ( .A1(n82), .A2(n53), .ZN(\ab[19][24] ) );
  NOR2_X1 U683 ( .A1(n175), .A2(n55), .ZN(\ab[17][26] ) );
  NOR2_X1 U684 ( .A1(n178), .A2(n57), .ZN(\ab[15][28] ) );
  NOR2_X1 U685 ( .A1(n136), .A2(n108), .ZN(\ab[3][14] ) );
  NOR2_X1 U686 ( .A1(n130), .A2(n112), .ZN(\ab[5][12] ) );
  NOR2_X1 U687 ( .A1(n124), .A2(n117), .ZN(\ab[7][10] ) );
  NOR2_X1 U688 ( .A1(n206), .A2(n200), .ZN(\ab[9][8] ) );
  NOR2_X1 U689 ( .A1(n196), .A2(n61), .ZN(\ab[11][6] ) );
  NOR2_X1 U690 ( .A1(n190), .A2(n59), .ZN(\ab[13][4] ) );
  NOR2_X1 U691 ( .A1(n183), .A2(n57), .ZN(\ab[15][2] ) );
  NOR2_X1 U692 ( .A1(n73), .A2(n51), .ZN(\ab[20][23] ) );
  NOR2_X1 U693 ( .A1(n172), .A2(n54), .ZN(\ab[18][25] ) );
  NOR2_X1 U694 ( .A1(n176), .A2(n56), .ZN(\ab[16][27] ) );
  NOR2_X1 U695 ( .A1(n133), .A2(n108), .ZN(\ab[3][13] ) );
  NOR2_X1 U696 ( .A1(n127), .A2(n112), .ZN(\ab[5][11] ) );
  NOR2_X1 U697 ( .A1(n203), .A2(n115), .ZN(\ab[7][9] ) );
  NOR2_X1 U698 ( .A1(n206), .A2(n197), .ZN(\ab[9][7] ) );
  NOR2_X1 U699 ( .A1(n193), .A2(n61), .ZN(\ab[11][5] ) );
  NOR2_X1 U700 ( .A1(n188), .A2(n59), .ZN(\ab[13][3] ) );
  NOR2_X1 U701 ( .A1(n156), .A2(n57), .ZN(\ab[15][1] ) );
  NOR2_X1 U702 ( .A1(n130), .A2(n108), .ZN(\ab[3][12] ) );
  NOR2_X1 U703 ( .A1(n124), .A2(n112), .ZN(\ab[5][10] ) );
  NOR2_X1 U704 ( .A1(n200), .A2(n115), .ZN(\ab[7][8] ) );
  NOR2_X1 U705 ( .A1(n206), .A2(n194), .ZN(\ab[9][6] ) );
  NOR2_X1 U706 ( .A1(n190), .A2(n61), .ZN(\ab[11][4] ) );
  NOR2_X1 U707 ( .A1(n183), .A2(n59), .ZN(\ab[13][2] ) );
  NOR2_X1 U708 ( .A1(n124), .A2(n110), .ZN(\ab[4][10] ) );
  NOR2_X1 U709 ( .A1(n200), .A2(n113), .ZN(\ab[6][8] ) );
  NOR2_X1 U710 ( .A1(n194), .A2(n118), .ZN(\ab[8][6] ) );
  NOR2_X1 U711 ( .A1(n190), .A2(n96), .ZN(\ab[10][4] ) );
  NOR2_X1 U712 ( .A1(n183), .A2(n60), .ZN(\ab[12][2] ) );
  NOR2_X1 U713 ( .A1(n163), .A2(n49), .ZN(\ab[22][22] ) );
  NOR2_X1 U714 ( .A1(n82), .A2(n51), .ZN(\ab[20][24] ) );
  NOR2_X1 U715 ( .A1(n173), .A2(n54), .ZN(\ab[18][26] ) );
  NOR2_X1 U716 ( .A1(n178), .A2(n56), .ZN(\ab[16][28] ) );
  NOR2_X1 U717 ( .A1(n124), .A2(n108), .ZN(\ab[3][10] ) );
  NOR2_X1 U718 ( .A1(n200), .A2(n111), .ZN(\ab[5][8] ) );
  NOR2_X1 U719 ( .A1(n194), .A2(n115), .ZN(\ab[7][6] ) );
  NOR2_X1 U720 ( .A1(n206), .A2(n189), .ZN(\ab[9][4] ) );
  NOR2_X1 U721 ( .A1(n183), .A2(n61), .ZN(\ab[11][2] ) );
  NOR2_X1 U722 ( .A1(n73), .A2(n50), .ZN(\ab[21][23] ) );
  NOR2_X1 U723 ( .A1(n170), .A2(n53), .ZN(\ab[19][25] ) );
  NOR2_X1 U724 ( .A1(n176), .A2(n55), .ZN(\ab[17][27] ) );
  NOR2_X1 U725 ( .A1(n203), .A2(n106), .ZN(\ab[3][9] ) );
  NOR2_X1 U726 ( .A1(n197), .A2(n111), .ZN(\ab[5][7] ) );
  NOR2_X1 U727 ( .A1(n191), .A2(n115), .ZN(\ab[7][5] ) );
  NOR2_X1 U728 ( .A1(n206), .A2(n186), .ZN(\ab[9][3] ) );
  NOR2_X1 U729 ( .A1(n156), .A2(n97), .ZN(\ab[11][1] ) );
  NOR2_X1 U730 ( .A1(n200), .A2(n106), .ZN(\ab[3][8] ) );
  NOR2_X1 U731 ( .A1(n194), .A2(n111), .ZN(\ab[5][6] ) );
  NOR2_X1 U732 ( .A1(n189), .A2(n115), .ZN(\ab[7][4] ) );
  NOR2_X1 U733 ( .A1(n206), .A2(n181), .ZN(\ab[9][2] ) );
  NOR2_X1 U734 ( .A1(n194), .A2(n109), .ZN(\ab[4][6] ) );
  NOR2_X1 U735 ( .A1(n189), .A2(n113), .ZN(\ab[6][4] ) );
  NOR2_X1 U736 ( .A1(n181), .A2(n118), .ZN(\ab[8][2] ) );
  NOR2_X1 U737 ( .A1(n194), .A2(n106), .ZN(\ab[3][6] ) );
  NOR2_X1 U738 ( .A1(n189), .A2(n111), .ZN(\ab[5][4] ) );
  NOR2_X1 U739 ( .A1(n181), .A2(n115), .ZN(\ab[7][2] ) );
  NOR2_X1 U740 ( .A1(n191), .A2(n106), .ZN(\ab[3][5] ) );
  NOR2_X1 U741 ( .A1(n186), .A2(n111), .ZN(\ab[5][3] ) );
  NOR2_X1 U742 ( .A1(n154), .A2(n116), .ZN(\ab[7][1] ) );
  NOR2_X1 U743 ( .A1(n167), .A2(n50), .ZN(\ab[21][24] ) );
  NOR2_X1 U744 ( .A1(n173), .A2(n53), .ZN(\ab[19][26] ) );
  NOR2_X1 U745 ( .A1(n177), .A2(n55), .ZN(\ab[17][28] ) );
  NOR2_X1 U746 ( .A1(n189), .A2(n106), .ZN(\ab[3][4] ) );
  NOR2_X1 U747 ( .A1(n181), .A2(n111), .ZN(\ab[5][2] ) );
  NOR2_X1 U748 ( .A1(n73), .A2(n49), .ZN(\ab[22][23] ) );
  NOR2_X1 U749 ( .A1(n170), .A2(n51), .ZN(\ab[20][25] ) );
  NOR2_X1 U750 ( .A1(n176), .A2(n54), .ZN(\ab[18][27] ) );
  NOR2_X1 U751 ( .A1(n186), .A2(n106), .ZN(\ab[3][3] ) );
  NOR2_X1 U752 ( .A1(n154), .A2(n112), .ZN(\ab[5][1] ) );
  NOR2_X1 U753 ( .A1(n181), .A2(n106), .ZN(\ab[3][2] ) );
  NOR2_X1 U754 ( .A1(n170), .A2(n50), .ZN(\ab[21][25] ) );
  NOR2_X1 U755 ( .A1(n176), .A2(n53), .ZN(\ab[19][27] ) );
  NOR2_X1 U756 ( .A1(n169), .A2(n49), .ZN(\ab[22][24] ) );
  NOR2_X1 U757 ( .A1(n175), .A2(n51), .ZN(\ab[20][26] ) );
  NOR2_X1 U758 ( .A1(n178), .A2(n54), .ZN(\ab[18][28] ) );
  NOR2_X1 U759 ( .A1(n189), .A2(n40), .ZN(\ab[30][4] ) );
  NOR2_X1 U760 ( .A1(n189), .A2(n42), .ZN(\ab[29][4] ) );
  NOR2_X1 U761 ( .A1(n191), .A2(n42), .ZN(\ab[29][5] ) );
  NOR2_X1 U762 ( .A1(n191), .A2(n43), .ZN(\ab[28][5] ) );
  NOR2_X1 U763 ( .A1(n200), .A2(n40), .ZN(\ab[30][8] ) );
  NOR2_X1 U764 ( .A1(n200), .A2(n42), .ZN(\ab[29][8] ) );
  NOR2_X1 U765 ( .A1(n203), .A2(n42), .ZN(\ab[29][9] ) );
  NOR2_X1 U766 ( .A1(n198), .A2(n45), .ZN(\ab[26][7] ) );
  NOR2_X1 U767 ( .A1(n186), .A2(n44), .ZN(\ab[27][3] ) );
  NOR2_X1 U768 ( .A1(n130), .A2(n42), .ZN(\ab[29][12] ) );
  NOR2_X1 U769 ( .A1(n154), .A2(n42), .ZN(\ab[29][1] ) );
  NOR2_X1 U770 ( .A1(n203), .A2(n43), .ZN(\ab[28][9] ) );
  NOR2_X1 U771 ( .A1(n121), .A2(n40), .ZN(\ab[30][0] ) );
  NOR2_X1 U772 ( .A1(n187), .A2(n45), .ZN(\ab[26][3] ) );
  NOR2_X1 U773 ( .A1(n127), .A2(n44), .ZN(\ab[27][11] ) );
  NOR2_X1 U774 ( .A1(n192), .A2(n47), .ZN(\ab[24][5] ) );
  NOR2_X1 U775 ( .A1(n154), .A2(n43), .ZN(\ab[28][1] ) );
  NOR2_X1 U776 ( .A1(n198), .A2(n48), .ZN(\ab[23][7] ) );
  NOR2_X1 U777 ( .A1(n128), .A2(n45), .ZN(\ab[26][11] ) );
  NOR2_X1 U778 ( .A1(n187), .A2(n46), .ZN(\ab[25][3] ) );
  NOR2_X1 U779 ( .A1(n198), .A2(n49), .ZN(\ab[22][7] ) );
  NOR2_X1 U780 ( .A1(n192), .A2(n48), .ZN(\ab[23][5] ) );
  NOR2_X1 U781 ( .A1(n121), .A2(n42), .ZN(\ab[29][0] ) );
  NOR2_X1 U782 ( .A1(n128), .A2(n48), .ZN(\ab[23][11] ) );
  NOR2_X1 U783 ( .A1(n204), .A2(n50), .ZN(\ab[21][9] ) );
  NOR2_X1 U784 ( .A1(n154), .A2(n44), .ZN(\ab[27][1] ) );
  NOR2_X1 U785 ( .A1(n198), .A2(n50), .ZN(\ab[21][7] ) );
  NOR2_X1 U786 ( .A1(n134), .A2(n47), .ZN(\ab[24][13] ) );
  NOR2_X1 U787 ( .A1(n128), .A2(n49), .ZN(\ab[22][11] ) );
  NOR2_X1 U788 ( .A1(n192), .A2(n49), .ZN(\ab[22][5] ) );
  NOR2_X1 U789 ( .A1(n187), .A2(n47), .ZN(\ab[24][3] ) );
  NOR2_X1 U790 ( .A1(n204), .A2(n51), .ZN(\ab[20][9] ) );
  NOR2_X1 U791 ( .A1(n140), .A2(n48), .ZN(\ab[23][15] ) );
  NOR2_X1 U792 ( .A1(n198), .A2(n51), .ZN(\ab[20][7] ) );
  NOR2_X1 U793 ( .A1(n204), .A2(n53), .ZN(\ab[19][9] ) );
  NOR2_X1 U794 ( .A1(n192), .A2(n50), .ZN(\ab[21][5] ) );
  NOR2_X1 U795 ( .A1(n128), .A2(n53), .ZN(\ab[19][11] ) );
  NOR2_X1 U796 ( .A1(n140), .A2(n49), .ZN(\ab[22][15] ) );
  NOR2_X1 U797 ( .A1(n121), .A2(n43), .ZN(\ab[28][0] ) );
  NOR2_X1 U798 ( .A1(n134), .A2(n50), .ZN(\ab[21][13] ) );
  NOR2_X1 U799 ( .A1(n155), .A2(n45), .ZN(\ab[26][1] ) );
  NOR2_X1 U800 ( .A1(n187), .A2(n48), .ZN(\ab[23][3] ) );
  NOR2_X1 U801 ( .A1(n198), .A2(n53), .ZN(\ab[19][7] ) );
  NOR2_X1 U802 ( .A1(n204), .A2(n54), .ZN(\ab[18][9] ) );
  NOR2_X1 U803 ( .A1(n128), .A2(n54), .ZN(\ab[18][11] ) );
  NOR2_X1 U804 ( .A1(n134), .A2(n51), .ZN(\ab[20][13] ) );
  NOR2_X1 U805 ( .A1(n146), .A2(n50), .ZN(\ab[21][17] ) );
  NOR2_X1 U806 ( .A1(n128), .A2(n55), .ZN(\ab[17][11] ) );
  NOR2_X1 U807 ( .A1(n192), .A2(n51), .ZN(\ab[20][5] ) );
  NOR2_X1 U808 ( .A1(n204), .A2(n55), .ZN(\ab[17][9] ) );
  NOR2_X1 U809 ( .A1(n198), .A2(n54), .ZN(\ab[18][7] ) );
  NOR2_X1 U810 ( .A1(n155), .A2(n46), .ZN(\ab[25][1] ) );
  NOR2_X1 U811 ( .A1(n187), .A2(n49), .ZN(\ab[22][3] ) );
  NOR2_X1 U812 ( .A1(n146), .A2(n51), .ZN(\ab[20][17] ) );
  NOR2_X1 U813 ( .A1(n128), .A2(n56), .ZN(\ab[16][11] ) );
  NOR2_X1 U814 ( .A1(n134), .A2(n55), .ZN(\ab[17][13] ) );
  NOR2_X1 U815 ( .A1(n140), .A2(n53), .ZN(\ab[19][15] ) );
  NOR2_X1 U816 ( .A1(n121), .A2(n44), .ZN(\ab[27][0] ) );
  NOR2_X1 U817 ( .A1(n204), .A2(n56), .ZN(\ab[16][9] ) );
  NOR2_X1 U818 ( .A1(n134), .A2(n56), .ZN(\ab[16][13] ) );
  NOR2_X1 U819 ( .A1(n195), .A2(n54), .ZN(\ab[18][6] ) );
  NOR2_X1 U820 ( .A1(n189), .A2(n51), .ZN(\ab[20][4] ) );
  NOR2_X1 U821 ( .A1(n140), .A2(n54), .ZN(\ab[18][15] ) );
  NOR2_X1 U822 ( .A1(n155), .A2(n47), .ZN(\ab[24][1] ) );
  NOR2_X1 U823 ( .A1(n129), .A2(n57), .ZN(\ab[15][11] ) );
  NOR2_X1 U824 ( .A1(n201), .A2(n56), .ZN(\ab[16][8] ) );
  NOR2_X1 U825 ( .A1(n135), .A2(n57), .ZN(\ab[15][13] ) );
  NOR2_X1 U826 ( .A1(n160), .A2(n119), .ZN(\ab[8][21] ) );
  NOR2_X1 U827 ( .A1(n207), .A2(n160), .ZN(\ab[9][21] ) );
  NOR2_X1 U828 ( .A1(n153), .A2(n96), .ZN(\ab[10][19] ) );
  NOR2_X1 U829 ( .A1(n153), .A2(n97), .ZN(\ab[11][19] ) );
  NOR2_X1 U830 ( .A1(n147), .A2(n98), .ZN(\ab[12][17] ) );
  NOR2_X1 U831 ( .A1(n147), .A2(n59), .ZN(\ab[13][17] ) );
  NOR2_X1 U832 ( .A1(n141), .A2(n99), .ZN(\ab[14][15] ) );
  NOR2_X1 U833 ( .A1(n141), .A2(n57), .ZN(\ab[15][15] ) );
  NOR2_X1 U834 ( .A1(n170), .A2(n119), .ZN(\ab[8][25] ) );
  NOR2_X1 U835 ( .A1(n207), .A2(n170), .ZN(\ab[9][25] ) );
  NOR2_X1 U836 ( .A1(n73), .A2(n97), .ZN(\ab[11][23] ) );
  NOR2_X1 U837 ( .A1(n162), .A2(n98), .ZN(\ab[12][21] ) );
  NOR2_X1 U838 ( .A1(n162), .A2(n59), .ZN(\ab[13][21] ) );
  NOR2_X1 U839 ( .A1(n153), .A2(n58), .ZN(\ab[14][19] ) );
  NOR2_X1 U840 ( .A1(n153), .A2(n57), .ZN(\ab[15][19] ) );
  NOR2_X1 U841 ( .A1(n146), .A2(n56), .ZN(\ab[16][17] ) );
  NOR2_X1 U842 ( .A1(n146), .A2(n55), .ZN(\ab[17][17] ) );
  NOR2_X1 U843 ( .A1(n170), .A2(n107), .ZN(\ab[3][25] ) );
  NOR2_X1 U844 ( .A1(n165), .A2(n112), .ZN(\ab[5][23] ) );
  NOR2_X1 U845 ( .A1(n160), .A2(n116), .ZN(\ab[7][21] ) );
  NOR2_X1 U846 ( .A1(n207), .A2(n151), .ZN(\ab[9][19] ) );
  NOR2_X1 U847 ( .A1(n147), .A2(n97), .ZN(\ab[11][17] ) );
  NOR2_X1 U848 ( .A1(n141), .A2(n59), .ZN(\ab[13][15] ) );
  NOR2_X1 U849 ( .A1(n182), .A2(n49), .ZN(\ab[22][2] ) );
  NOR2_X1 U850 ( .A1(n160), .A2(n114), .ZN(\ab[6][21] ) );
  NOR2_X1 U851 ( .A1(n151), .A2(n119), .ZN(\ab[8][19] ) );
  NOR2_X1 U852 ( .A1(n147), .A2(n62), .ZN(\ab[10][17] ) );
  NOR2_X1 U853 ( .A1(n141), .A2(n98), .ZN(\ab[12][15] ) );
  NOR2_X1 U854 ( .A1(n135), .A2(n99), .ZN(\ab[14][13] ) );
  NOR2_X1 U855 ( .A1(n152), .A2(n54), .ZN(\ab[18][19] ) );
  NOR2_X1 U856 ( .A1(n165), .A2(n107), .ZN(\ab[3][23] ) );
  NOR2_X1 U857 ( .A1(n160), .A2(n112), .ZN(\ab[5][21] ) );
  NOR2_X1 U858 ( .A1(n151), .A2(n116), .ZN(\ab[7][19] ) );
  NOR2_X1 U859 ( .A1(n207), .A2(n145), .ZN(\ab[9][17] ) );
  NOR2_X1 U860 ( .A1(n141), .A2(n97), .ZN(\ab[11][15] ) );
  NOR2_X1 U861 ( .A1(n135), .A2(n59), .ZN(\ab[13][13] ) );
  NOR2_X1 U862 ( .A1(n160), .A2(n110), .ZN(\ab[4][21] ) );
  NOR2_X1 U863 ( .A1(n151), .A2(n114), .ZN(\ab[6][19] ) );
  NOR2_X1 U864 ( .A1(n145), .A2(n119), .ZN(\ab[8][17] ) );
  NOR2_X1 U865 ( .A1(n141), .A2(n96), .ZN(\ab[10][15] ) );
  NOR2_X1 U866 ( .A1(n135), .A2(n98), .ZN(\ab[12][13] ) );
  NOR2_X1 U867 ( .A1(n129), .A2(n99), .ZN(\ab[14][11] ) );
  NOR2_X1 U868 ( .A1(n157), .A2(n110), .ZN(\ab[4][20] ) );
  NOR2_X1 U869 ( .A1(n148), .A2(n114), .ZN(\ab[6][18] ) );
  NOR2_X1 U870 ( .A1(n142), .A2(n119), .ZN(\ab[8][16] ) );
  NOR2_X1 U871 ( .A1(n138), .A2(n96), .ZN(\ab[10][14] ) );
  NOR2_X1 U872 ( .A1(n132), .A2(n60), .ZN(\ab[12][12] ) );
  NOR2_X1 U873 ( .A1(n126), .A2(n99), .ZN(\ab[14][10] ) );
  NOR2_X1 U874 ( .A1(n151), .A2(n110), .ZN(\ab[4][19] ) );
  NOR2_X1 U875 ( .A1(n145), .A2(n114), .ZN(\ab[6][17] ) );
  NOR2_X1 U876 ( .A1(n139), .A2(n120), .ZN(\ab[8][15] ) );
  NOR2_X1 U877 ( .A1(n135), .A2(n96), .ZN(\ab[10][13] ) );
  NOR2_X1 U878 ( .A1(n129), .A2(n60), .ZN(\ab[12][11] ) );
  NOR2_X1 U879 ( .A1(n205), .A2(n58), .ZN(\ab[14][9] ) );
  NOR2_X1 U880 ( .A1(n198), .A2(n56), .ZN(\ab[16][7] ) );
  NOR2_X1 U881 ( .A1(n192), .A2(n54), .ZN(\ab[18][5] ) );
  NOR2_X1 U882 ( .A1(n187), .A2(n51), .ZN(\ab[20][3] ) );
  NOR2_X1 U883 ( .A1(n155), .A2(n49), .ZN(\ab[22][1] ) );
  NOR2_X1 U884 ( .A1(n148), .A2(n110), .ZN(\ab[4][18] ) );
  NOR2_X1 U885 ( .A1(n142), .A2(n114), .ZN(\ab[6][16] ) );
  NOR2_X1 U886 ( .A1(n136), .A2(n120), .ZN(\ab[8][14] ) );
  NOR2_X1 U887 ( .A1(n132), .A2(n96), .ZN(\ab[10][12] ) );
  NOR2_X1 U888 ( .A1(n126), .A2(n60), .ZN(\ab[12][10] ) );
  NOR2_X1 U889 ( .A1(n202), .A2(n58), .ZN(\ab[14][8] ) );
  NOR2_X1 U890 ( .A1(n195), .A2(n56), .ZN(\ab[16][6] ) );
  NOR2_X1 U891 ( .A1(n189), .A2(n54), .ZN(\ab[18][4] ) );
  NOR2_X1 U892 ( .A1(n182), .A2(n51), .ZN(\ab[20][2] ) );
  NOR2_X1 U893 ( .A1(n151), .A2(n105), .ZN(\ab[2][19] ) );
  AND2_X1 U894 ( .A1(\ab[1][19] ), .A2(\ab[0][20] ), .ZN(\CARRYB[1][19] ) );
  NOR2_X1 U895 ( .A1(n145), .A2(n110), .ZN(\ab[4][17] ) );
  NOR2_X1 U896 ( .A1(n139), .A2(n114), .ZN(\ab[6][15] ) );
  NOR2_X1 U897 ( .A1(n133), .A2(n120), .ZN(\ab[8][13] ) );
  NOR2_X1 U898 ( .A1(n129), .A2(n96), .ZN(\ab[10][11] ) );
  NOR2_X1 U899 ( .A1(n205), .A2(n60), .ZN(\ab[12][9] ) );
  NOR2_X1 U900 ( .A1(n199), .A2(n58), .ZN(\ab[14][7] ) );
  NOR2_X1 U901 ( .A1(n192), .A2(n56), .ZN(\ab[16][5] ) );
  NOR2_X1 U902 ( .A1(n187), .A2(n54), .ZN(\ab[18][3] ) );
  NOR2_X1 U903 ( .A1(n155), .A2(n51), .ZN(\ab[20][1] ) );
  NOR2_X1 U904 ( .A1(n148), .A2(n104), .ZN(\ab[2][18] ) );
  AND2_X1 U905 ( .A1(\ab[1][18] ), .A2(\ab[0][19] ), .ZN(\CARRYB[1][18] ) );
  NOR2_X1 U906 ( .A1(n142), .A2(n110), .ZN(\ab[4][16] ) );
  NOR2_X1 U907 ( .A1(n136), .A2(n114), .ZN(\ab[6][14] ) );
  NOR2_X1 U908 ( .A1(n130), .A2(n120), .ZN(\ab[8][12] ) );
  NOR2_X1 U909 ( .A1(n126), .A2(n96), .ZN(\ab[10][10] ) );
  NOR2_X1 U910 ( .A1(n202), .A2(n60), .ZN(\ab[12][8] ) );
  NOR2_X1 U911 ( .A1(n196), .A2(n58), .ZN(\ab[14][6] ) );
  NOR2_X1 U912 ( .A1(n189), .A2(n56), .ZN(\ab[16][4] ) );
  NOR2_X1 U913 ( .A1(n182), .A2(n54), .ZN(\ab[18][2] ) );
  NOR2_X1 U914 ( .A1(n145), .A2(n104), .ZN(\ab[2][17] ) );
  AND2_X1 U915 ( .A1(\ab[1][17] ), .A2(\ab[0][18] ), .ZN(\CARRYB[1][17] ) );
  NOR2_X1 U916 ( .A1(n139), .A2(n110), .ZN(\ab[4][15] ) );
  NOR2_X1 U917 ( .A1(n133), .A2(n114), .ZN(\ab[6][13] ) );
  NOR2_X1 U918 ( .A1(n127), .A2(n120), .ZN(\ab[8][11] ) );
  NOR2_X1 U919 ( .A1(n205), .A2(n96), .ZN(\ab[10][9] ) );
  NOR2_X1 U920 ( .A1(n199), .A2(n60), .ZN(\ab[12][7] ) );
  NOR2_X1 U921 ( .A1(n193), .A2(n58), .ZN(\ab[14][5] ) );
  NOR2_X1 U922 ( .A1(n187), .A2(n56), .ZN(\ab[16][3] ) );
  NOR2_X1 U923 ( .A1(n155), .A2(n54), .ZN(\ab[18][1] ) );
  NOR2_X1 U924 ( .A1(n142), .A2(n105), .ZN(\ab[2][16] ) );
  AND2_X1 U925 ( .A1(\ab[1][16] ), .A2(\ab[0][17] ), .ZN(\CARRYB[1][16] ) );
  NOR2_X1 U926 ( .A1(n136), .A2(n110), .ZN(\ab[4][14] ) );
  NOR2_X1 U927 ( .A1(n130), .A2(n114), .ZN(\ab[6][12] ) );
  NOR2_X1 U928 ( .A1(n124), .A2(n120), .ZN(\ab[8][10] ) );
  NOR2_X1 U929 ( .A1(n202), .A2(n96), .ZN(\ab[10][8] ) );
  NOR2_X1 U930 ( .A1(n196), .A2(n60), .ZN(\ab[12][6] ) );
  NOR2_X1 U931 ( .A1(n190), .A2(n58), .ZN(\ab[14][4] ) );
  NOR2_X1 U932 ( .A1(n182), .A2(n56), .ZN(\ab[16][2] ) );
  NOR2_X1 U933 ( .A1(n139), .A2(n104), .ZN(\ab[2][15] ) );
  AND2_X1 U934 ( .A1(\ab[1][15] ), .A2(\ab[0][16] ), .ZN(\CARRYB[1][15] ) );
  NOR2_X1 U935 ( .A1(n133), .A2(n110), .ZN(\ab[4][13] ) );
  NOR2_X1 U936 ( .A1(n127), .A2(n114), .ZN(\ab[6][11] ) );
  NOR2_X1 U937 ( .A1(n203), .A2(n118), .ZN(\ab[8][9] ) );
  NOR2_X1 U938 ( .A1(n199), .A2(n96), .ZN(\ab[10][7] ) );
  NOR2_X1 U939 ( .A1(n193), .A2(n60), .ZN(\ab[12][5] ) );
  NOR2_X1 U940 ( .A1(n188), .A2(n58), .ZN(\ab[14][3] ) );
  NOR2_X1 U941 ( .A1(n155), .A2(n56), .ZN(\ab[16][1] ) );
  NOR2_X1 U942 ( .A1(n136), .A2(n104), .ZN(\ab[2][14] ) );
  AND2_X1 U943 ( .A1(\ab[1][14] ), .A2(\ab[0][15] ), .ZN(\CARRYB[1][14] ) );
  NOR2_X1 U944 ( .A1(n130), .A2(n110), .ZN(\ab[4][12] ) );
  NOR2_X1 U945 ( .A1(n124), .A2(n114), .ZN(\ab[6][10] ) );
  NOR2_X1 U946 ( .A1(n200), .A2(n118), .ZN(\ab[8][8] ) );
  NOR2_X1 U947 ( .A1(n196), .A2(n96), .ZN(\ab[10][6] ) );
  NOR2_X1 U948 ( .A1(n190), .A2(n60), .ZN(\ab[12][4] ) );
  NOR2_X1 U949 ( .A1(n183), .A2(n58), .ZN(\ab[14][2] ) );
  NOR2_X1 U950 ( .A1(n133), .A2(n105), .ZN(\ab[2][13] ) );
  AND2_X1 U951 ( .A1(\ab[1][13] ), .A2(\ab[0][14] ), .ZN(\CARRYB[1][13] ) );
  NOR2_X1 U952 ( .A1(n127), .A2(n110), .ZN(\ab[4][11] ) );
  NOR2_X1 U953 ( .A1(n203), .A2(n113), .ZN(\ab[6][9] ) );
  NOR2_X1 U954 ( .A1(n197), .A2(n118), .ZN(\ab[8][7] ) );
  NOR2_X1 U955 ( .A1(n193), .A2(n96), .ZN(\ab[10][5] ) );
  NOR2_X1 U956 ( .A1(n188), .A2(n60), .ZN(\ab[12][3] ) );
  NOR2_X1 U957 ( .A1(n156), .A2(n58), .ZN(\ab[14][1] ) );
  NOR2_X1 U958 ( .A1(n127), .A2(n108), .ZN(\ab[3][11] ) );
  NOR2_X1 U959 ( .A1(n127), .A2(n105), .ZN(\ab[2][11] ) );
  AND2_X1 U960 ( .A1(\ab[1][11] ), .A2(\ab[0][12] ), .ZN(\CARRYB[1][11] ) );
  NOR2_X1 U961 ( .A1(n203), .A2(n111), .ZN(\ab[5][9] ) );
  NOR2_X1 U962 ( .A1(n203), .A2(n109), .ZN(\ab[4][9] ) );
  NOR2_X1 U963 ( .A1(n197), .A2(n115), .ZN(\ab[7][7] ) );
  NOR2_X1 U964 ( .A1(n197), .A2(n113), .ZN(\ab[6][7] ) );
  NOR2_X1 U965 ( .A1(n206), .A2(n191), .ZN(\ab[9][5] ) );
  NOR2_X1 U966 ( .A1(n191), .A2(n118), .ZN(\ab[8][5] ) );
  NOR2_X1 U967 ( .A1(n188), .A2(n61), .ZN(\ab[11][3] ) );
  NOR2_X1 U968 ( .A1(n188), .A2(n96), .ZN(\ab[10][3] ) );
  NOR2_X1 U969 ( .A1(n156), .A2(n59), .ZN(\ab[13][1] ) );
  NOR2_X1 U970 ( .A1(n130), .A2(n104), .ZN(\ab[2][12] ) );
  AND2_X1 U971 ( .A1(\ab[1][12] ), .A2(\ab[0][13] ), .ZN(\CARRYB[1][12] ) );
  NOR2_X1 U972 ( .A1(n156), .A2(n98), .ZN(\ab[12][1] ) );
  NOR2_X1 U973 ( .A1(n124), .A2(n105), .ZN(\ab[2][10] ) );
  AND2_X1 U974 ( .A1(\ab[1][10] ), .A2(\ab[0][11] ), .ZN(\CARRYB[1][10] ) );
  NOR2_X1 U975 ( .A1(n200), .A2(n109), .ZN(\ab[4][8] ) );
  NOR2_X1 U976 ( .A1(n194), .A2(n113), .ZN(\ab[6][6] ) );
  NOR2_X1 U977 ( .A1(n189), .A2(n118), .ZN(\ab[8][4] ) );
  NOR2_X1 U978 ( .A1(n183), .A2(n96), .ZN(\ab[10][2] ) );
  NOR2_X1 U979 ( .A1(n203), .A2(n104), .ZN(\ab[2][9] ) );
  AND2_X1 U980 ( .A1(\ab[1][9] ), .A2(\ab[0][10] ), .ZN(\CARRYB[1][9] ) );
  NOR2_X1 U981 ( .A1(n197), .A2(n109), .ZN(\ab[4][7] ) );
  NOR2_X1 U982 ( .A1(n191), .A2(n113), .ZN(\ab[6][5] ) );
  NOR2_X1 U983 ( .A1(n186), .A2(n118), .ZN(\ab[8][3] ) );
  NOR2_X1 U984 ( .A1(n156), .A2(n62), .ZN(\ab[10][1] ) );
  NOR2_X1 U985 ( .A1(n197), .A2(n106), .ZN(\ab[3][7] ) );
  NOR2_X1 U986 ( .A1(n197), .A2(n104), .ZN(\ab[2][7] ) );
  AND2_X1 U987 ( .A1(\ab[1][7] ), .A2(\ab[0][8] ), .ZN(\CARRYB[1][7] ) );
  NOR2_X1 U988 ( .A1(n191), .A2(n111), .ZN(\ab[5][5] ) );
  NOR2_X1 U989 ( .A1(n191), .A2(n109), .ZN(\ab[4][5] ) );
  NOR2_X1 U990 ( .A1(n186), .A2(n115), .ZN(\ab[7][3] ) );
  NOR2_X1 U991 ( .A1(n186), .A2(n113), .ZN(\ab[6][3] ) );
  NOR2_X1 U992 ( .A1(n207), .A2(n154), .ZN(\ab[9][1] ) );
  NOR2_X1 U993 ( .A1(n154), .A2(n119), .ZN(\ab[8][1] ) );
  NOR2_X1 U994 ( .A1(n194), .A2(n104), .ZN(\ab[2][6] ) );
  AND2_X1 U995 ( .A1(\ab[1][6] ), .A2(\ab[0][7] ), .ZN(\CARRYB[1][6] ) );
  NOR2_X1 U996 ( .A1(n189), .A2(n109), .ZN(\ab[4][4] ) );
  NOR2_X1 U997 ( .A1(n181), .A2(n113), .ZN(\ab[6][2] ) );
  NOR2_X1 U998 ( .A1(n191), .A2(n105), .ZN(\ab[2][5] ) );
  AND2_X1 U999 ( .A1(\ab[1][5] ), .A2(\ab[0][6] ), .ZN(\CARRYB[1][5] ) );
  NOR2_X1 U1000 ( .A1(n186), .A2(n109), .ZN(\ab[4][3] ) );
  NOR2_X1 U1001 ( .A1(n154), .A2(n114), .ZN(\ab[6][1] ) );
  NOR2_X1 U1002 ( .A1(n189), .A2(n104), .ZN(\ab[2][4] ) );
  AND2_X1 U1003 ( .A1(\ab[1][4] ), .A2(\ab[0][5] ), .ZN(\CARRYB[1][4] ) );
  NOR2_X1 U1004 ( .A1(n181), .A2(n109), .ZN(\ab[4][2] ) );
  NOR2_X1 U1005 ( .A1(n186), .A2(n105), .ZN(\ab[2][3] ) );
  AND2_X1 U1006 ( .A1(\ab[1][3] ), .A2(\ab[0][4] ), .ZN(\CARRYB[1][3] ) );
  NOR2_X1 U1007 ( .A1(n154), .A2(n110), .ZN(\ab[4][1] ) );
  NOR2_X1 U1008 ( .A1(n154), .A2(n107), .ZN(\ab[3][1] ) );
  NOR2_X1 U1009 ( .A1(n154), .A2(n105), .ZN(\ab[2][1] ) );
  AND2_X1 U1010 ( .A1(\ab[1][1] ), .A2(\ab[0][2] ), .ZN(\CARRYB[1][1] ) );
  NOR2_X1 U1011 ( .A1(n122), .A2(n45), .ZN(\ab[26][0] ) );
  NOR2_X1 U1012 ( .A1(n122), .A2(n46), .ZN(\ab[25][0] ) );
  NOR2_X1 U1013 ( .A1(n122), .A2(n47), .ZN(\ab[24][0] ) );
  NOR2_X1 U1014 ( .A1(n122), .A2(n48), .ZN(\ab[23][0] ) );
  NOR2_X1 U1015 ( .A1(n122), .A2(n49), .ZN(\ab[22][0] ) );
  NOR2_X1 U1016 ( .A1(n122), .A2(n50), .ZN(\ab[21][0] ) );
  NOR2_X1 U1017 ( .A1(n122), .A2(n51), .ZN(\ab[20][0] ) );
  NOR2_X1 U1018 ( .A1(n122), .A2(n53), .ZN(\ab[19][0] ) );
  NOR2_X1 U1019 ( .A1(n122), .A2(n54), .ZN(\ab[18][0] ) );
  NOR2_X1 U1020 ( .A1(n122), .A2(n55), .ZN(\ab[17][0] ) );
  NOR2_X1 U1021 ( .A1(n122), .A2(n56), .ZN(\ab[16][0] ) );
  NOR2_X1 U1022 ( .A1(n123), .A2(n57), .ZN(\ab[15][0] ) );
  NOR2_X1 U1023 ( .A1(n123), .A2(n99), .ZN(\ab[14][0] ) );
  NOR2_X1 U1024 ( .A1(n123), .A2(n59), .ZN(\ab[13][0] ) );
  NOR2_X1 U1025 ( .A1(n123), .A2(n60), .ZN(\ab[12][0] ) );
  NOR2_X1 U1026 ( .A1(n123), .A2(n61), .ZN(\ab[11][0] ) );
  NOR2_X1 U1027 ( .A1(n123), .A2(n96), .ZN(\ab[10][0] ) );
  NOR2_X1 U1028 ( .A1(n2), .A2(n121), .ZN(\ab[9][0] ) );
  NOR2_X1 U1029 ( .A1(n121), .A2(n120), .ZN(\ab[8][0] ) );
  NOR2_X1 U1030 ( .A1(n121), .A2(n117), .ZN(\ab[7][0] ) );
  NOR2_X1 U1031 ( .A1(n121), .A2(n114), .ZN(\ab[6][0] ) );
  NOR2_X1 U1032 ( .A1(n121), .A2(n112), .ZN(\ab[5][0] ) );
  NOR2_X1 U1033 ( .A1(n121), .A2(n110), .ZN(\ab[4][0] ) );
  NOR2_X1 U1034 ( .A1(n121), .A2(n108), .ZN(\ab[3][0] ) );
  NOR2_X1 U1035 ( .A1(n121), .A2(n104), .ZN(\ab[2][0] ) );
  AND2_X1 U1036 ( .A1(\ab[1][0] ), .A2(\ab[0][1] ), .ZN(\CARRYB[1][0] ) );
  NOR2_X1 U1037 ( .A1(n181), .A2(n104), .ZN(\ab[2][2] ) );
  AND2_X1 U1038 ( .A1(\ab[1][2] ), .A2(\ab[0][3] ), .ZN(\CARRYB[1][2] ) );
  NOR2_X1 U1039 ( .A1(n160), .A2(n40), .ZN(\ab[30][21] ) );
  NOR2_X1 U1040 ( .A1(n164), .A2(n40), .ZN(\ab[30][22] ) );
  NOR2_X1 U1041 ( .A1(n157), .A2(n40), .ZN(\ab[30][20] ) );
  NOR2_X1 U1042 ( .A1(n165), .A2(n40), .ZN(\ab[30][23] ) );
  NOR2_X1 U1043 ( .A1(n151), .A2(n40), .ZN(\ab[30][19] ) );
  NOR2_X1 U1044 ( .A1(n160), .A2(n42), .ZN(\ab[29][21] ) );
  NOR2_X1 U1045 ( .A1(n164), .A2(n42), .ZN(\ab[29][22] ) );
  NOR2_X1 U1046 ( .A1(n157), .A2(n42), .ZN(\ab[29][20] ) );
  NOR2_X1 U1047 ( .A1(n165), .A2(n42), .ZN(\ab[29][23] ) );
  NOR2_X1 U1048 ( .A1(n169), .A2(n40), .ZN(\ab[30][24] ) );
  NOR2_X1 U1049 ( .A1(n148), .A2(n40), .ZN(\ab[30][18] ) );
  NOR2_X1 U1050 ( .A1(n163), .A2(n43), .ZN(\ab[28][22] ) );
  NOR2_X1 U1051 ( .A1(n160), .A2(n43), .ZN(\ab[28][21] ) );
  NOR2_X1 U1052 ( .A1(n151), .A2(n42), .ZN(\ab[29][19] ) );
  NOR2_X1 U1053 ( .A1(n167), .A2(n42), .ZN(\ab[29][24] ) );
  NOR2_X1 U1054 ( .A1(n165), .A2(n43), .ZN(\ab[28][23] ) );
  NOR2_X1 U1055 ( .A1(n157), .A2(n43), .ZN(\ab[28][20] ) );
  NOR2_X1 U1056 ( .A1(n82), .A2(n43), .ZN(\ab[28][24] ) );
  NOR2_X1 U1057 ( .A1(n163), .A2(n44), .ZN(\ab[27][22] ) );
  NOR2_X1 U1058 ( .A1(n160), .A2(n44), .ZN(\ab[27][21] ) );
  NOR2_X1 U1059 ( .A1(n165), .A2(n44), .ZN(\ab[27][23] ) );
  NOR2_X1 U1060 ( .A1(n172), .A2(n40), .ZN(\ab[30][25] ) );
  NOR2_X1 U1061 ( .A1(n151), .A2(n43), .ZN(\ab[28][19] ) );
  NOR2_X1 U1062 ( .A1(n148), .A2(n42), .ZN(\ab[29][18] ) );
  NOR2_X1 U1063 ( .A1(n170), .A2(n42), .ZN(\ab[29][25] ) );
  NOR2_X1 U1064 ( .A1(n82), .A2(n44), .ZN(\ab[27][24] ) );
  NOR2_X1 U1065 ( .A1(n157), .A2(n44), .ZN(\ab[27][20] ) );
  NOR2_X1 U1066 ( .A1(n164), .A2(n45), .ZN(\ab[26][22] ) );
  NOR2_X1 U1067 ( .A1(n73), .A2(n45), .ZN(\ab[26][23] ) );
  NOR2_X1 U1068 ( .A1(n172), .A2(n43), .ZN(\ab[28][25] ) );
  NOR2_X1 U1069 ( .A1(n145), .A2(n40), .ZN(\ab[30][17] ) );
  NOR2_X1 U1070 ( .A1(n161), .A2(n45), .ZN(\ab[26][21] ) );
  NOR2_X1 U1071 ( .A1(n169), .A2(n45), .ZN(\ab[26][24] ) );
  NOR2_X1 U1072 ( .A1(n170), .A2(n44), .ZN(\ab[27][25] ) );
  NOR2_X1 U1073 ( .A1(n175), .A2(n40), .ZN(\ab[30][26] ) );
  NOR2_X1 U1074 ( .A1(n73), .A2(n46), .ZN(\ab[25][23] ) );
  NOR2_X1 U1075 ( .A1(n163), .A2(n46), .ZN(\ab[25][22] ) );
  NOR2_X1 U1076 ( .A1(n176), .A2(n40), .ZN(\ab[30][27] ) );
  NOR2_X1 U1077 ( .A1(n170), .A2(n45), .ZN(\ab[26][25] ) );
  NOR2_X1 U1078 ( .A1(n167), .A2(n46), .ZN(\ab[25][24] ) );
  NOR2_X1 U1079 ( .A1(n177), .A2(n40), .ZN(\ab[30][28] ) );
  NOR2_X1 U1080 ( .A1(n173), .A2(n42), .ZN(\ab[29][26] ) );
  NOR2_X1 U1081 ( .A1(n175), .A2(n43), .ZN(\ab[28][26] ) );
  NOR2_X1 U1082 ( .A1(n73), .A2(n47), .ZN(\ab[24][23] ) );
  NOR2_X1 U1083 ( .A1(n170), .A2(n46), .ZN(\ab[25][25] ) );
  NOR2_X1 U1084 ( .A1(n82), .A2(n47), .ZN(\ab[24][24] ) );
  NOR2_X1 U1085 ( .A1(n173), .A2(n44), .ZN(\ab[27][26] ) );
  NOR2_X1 U1086 ( .A1(n173), .A2(n45), .ZN(\ab[26][26] ) );
  NOR2_X1 U1087 ( .A1(n170), .A2(n47), .ZN(\ab[24][25] ) );
  NOR2_X1 U1088 ( .A1(n82), .A2(n48), .ZN(\ab[23][24] ) );
  NOR2_X1 U1089 ( .A1(n176), .A2(n42), .ZN(\ab[29][27] ) );
  NOR2_X1 U1090 ( .A1(n175), .A2(n46), .ZN(\ab[25][26] ) );
  NOR2_X1 U1091 ( .A1(n172), .A2(n48), .ZN(\ab[23][25] ) );
  NOR2_X1 U1092 ( .A1(n173), .A2(n47), .ZN(\ab[24][26] ) );
  NOR2_X1 U1093 ( .A1(n177), .A2(n42), .ZN(\ab[29][28] ) );
  NOR2_X1 U1094 ( .A1(n173), .A2(n50), .ZN(\ab[21][26] ) );
  NOR2_X1 U1095 ( .A1(n178), .A2(n53), .ZN(\ab[19][28] ) );
  NOR2_X1 U1096 ( .A1(n170), .A2(n49), .ZN(\ab[22][25] ) );
  NOR2_X1 U1097 ( .A1(n176), .A2(n51), .ZN(\ab[20][27] ) );
  NOR2_X1 U1098 ( .A1(n176), .A2(n43), .ZN(\ab[28][27] ) );
  NOR2_X1 U1099 ( .A1(n176), .A2(n50), .ZN(\ab[21][27] ) );
  NOR2_X1 U1100 ( .A1(n175), .A2(n49), .ZN(\ab[22][26] ) );
  NOR2_X1 U1101 ( .A1(n177), .A2(n51), .ZN(\ab[20][28] ) );
  NOR2_X1 U1102 ( .A1(n173), .A2(n48), .ZN(\ab[23][26] ) );
  NOR2_X1 U1103 ( .A1(n176), .A2(n44), .ZN(\ab[27][27] ) );
  NOR2_X1 U1104 ( .A1(n176), .A2(n45), .ZN(\ab[26][27] ) );
  NOR2_X1 U1105 ( .A1(n178), .A2(n50), .ZN(\ab[21][28] ) );
  NOR2_X1 U1106 ( .A1(n176), .A2(n49), .ZN(\ab[22][27] ) );
  NOR2_X1 U1107 ( .A1(n176), .A2(n46), .ZN(\ab[25][27] ) );
  NOR2_X1 U1108 ( .A1(n176), .A2(n48), .ZN(\ab[23][27] ) );
  NOR2_X1 U1109 ( .A1(n178), .A2(n49), .ZN(\ab[22][28] ) );
  NOR2_X1 U1110 ( .A1(n176), .A2(n47), .ZN(\ab[24][27] ) );
  NOR2_X1 U1111 ( .A1(n177), .A2(n48), .ZN(\ab[23][28] ) );
  NOR2_X1 U1112 ( .A1(n178), .A2(n47), .ZN(\ab[24][28] ) );
  NOR2_X1 U1113 ( .A1(n178), .A2(n46), .ZN(\ab[25][28] ) );
  NOR2_X1 U1114 ( .A1(n177), .A2(n45), .ZN(\ab[26][28] ) );
  NOR2_X1 U1115 ( .A1(n178), .A2(n43), .ZN(\ab[28][28] ) );
  NOR2_X1 U1116 ( .A1(n178), .A2(n44), .ZN(\ab[27][28] ) );
  NOR2_X1 U1117 ( .A1(n209), .A2(QA), .ZN(\ab[31][31] ) );
  NOR2_X1 U1118 ( .A1(n123), .A2(n94), .ZN(PRODUCT[0]) );
  CLKBUF_X3 U1119 ( .A(n7), .Z(n191) );
  CLKBUF_X3 U1120 ( .A(n6), .Z(n194) );
  CLKBUF_X3 U1121 ( .A(n9), .Z(n186) );
  CLKBUF_X3 U1122 ( .A(n19), .Z(n163) );
  CLKBUF_X3 U1123 ( .A(n20), .Z(n160) );
  CLKBUF_X3 U1124 ( .A(n5), .Z(n197) );
  CLKBUF_X3 U1125 ( .A(n28), .Z(n136) );
  CLKBUF_X3 U1126 ( .A(n11), .Z(n181) );
  CLKBUF_X3 U1127 ( .A(n27), .Z(n139) );
  CLKBUF_X3 U1128 ( .A(n18), .Z(n165) );
  CLKBUF_X3 U1129 ( .A(n21), .Z(n157) );
  CLKBUF_X3 U1130 ( .A(n4), .Z(n200) );
  CLKBUF_X3 U1131 ( .A(n29), .Z(n133) );
  CLKBUF_X3 U1132 ( .A(n3), .Z(n203) );
  CLKBUF_X3 U1133 ( .A(n32), .Z(n124) );
  CLKBUF_X3 U1134 ( .A(n30), .Z(n130) );
  CLKBUF_X3 U1135 ( .A(n31), .Z(n127) );
  CLKBUF_X3 U1136 ( .A(n26), .Z(n142) );
  CLKBUF_X3 U1137 ( .A(n23), .Z(n151) );
  CLKBUF_X3 U1138 ( .A(n6), .Z(n195) );
  CLKBUF_X3 U1139 ( .A(n4), .Z(n201) );
  CLKBUF_X3 U1140 ( .A(n7), .Z(n192) );
  BUF_X2 U1141 ( .A(n23), .Z(n152) );
  BUF_X2 U1142 ( .A(n11), .Z(n182) );
  CLKBUF_X1 U1143 ( .A(n39), .Z(n108) );
  BUF_X1 U1144 ( .A(n20), .Z(n162) );
  BUF_X1 U1145 ( .A(n21), .Z(n159) );
  BUF_X1 U1146 ( .A(n23), .Z(n153) );
  BUF_X1 U1147 ( .A(n24), .Z(n150) );
  BUF_X1 U1148 ( .A(n25), .Z(n147) );
  BUF_X1 U1149 ( .A(n26), .Z(n144) );
  BUF_X1 U1150 ( .A(n27), .Z(n141) );
  BUF_X1 U1151 ( .A(n29), .Z(n135) );
  BUF_X1 U1152 ( .A(n28), .Z(n138) );
  BUF_X1 U1153 ( .A(n30), .Z(n132) );
  BUF_X1 U1154 ( .A(n31), .Z(n129) );
  BUF_X1 U1155 ( .A(n32), .Z(n126) );
  BUF_X1 U1156 ( .A(n3), .Z(n205) );
  BUF_X1 U1157 ( .A(n4), .Z(n202) );
  BUF_X1 U1158 ( .A(n5), .Z(n199) );
  BUF_X1 U1159 ( .A(n6), .Z(n196) );
  BUF_X1 U1160 ( .A(n7), .Z(n193) );
  BUF_X1 U1161 ( .A(n8), .Z(n190) );
  BUF_X1 U1162 ( .A(n11), .Z(n183) );
  BUF_X1 U1163 ( .A(n9), .Z(n188) );
  BUF_X1 U1164 ( .A(n22), .Z(n156) );
  AND2_X1 U1165 ( .A1(\ab[1][29] ), .A2(\ab[0][30] ), .ZN(\CARRYB[1][29] ) );
  NOR2_X1 U1166 ( .A1(n180), .A2(n106), .ZN(\ab[3][29] ) );
  NOR2_X1 U1167 ( .A1(n180), .A2(n109), .ZN(\ab[4][29] ) );
  NOR2_X1 U1168 ( .A1(n180), .A2(n111), .ZN(\ab[5][29] ) );
  NOR2_X1 U1169 ( .A1(n180), .A2(n113), .ZN(\ab[6][29] ) );
  NOR2_X1 U1170 ( .A1(n180), .A2(n115), .ZN(\ab[7][29] ) );
  NOR2_X1 U1171 ( .A1(n180), .A2(n118), .ZN(\ab[8][29] ) );
  NOR2_X1 U1172 ( .A1(n206), .A2(n180), .ZN(\ab[9][29] ) );
  NOR2_X1 U1173 ( .A1(n180), .A2(n62), .ZN(\ab[10][29] ) );
  NOR2_X1 U1174 ( .A1(n180), .A2(n61), .ZN(\ab[11][29] ) );
  NOR2_X1 U1175 ( .A1(n180), .A2(n60), .ZN(\ab[12][29] ) );
  NOR2_X1 U1176 ( .A1(n180), .A2(n59), .ZN(\ab[13][29] ) );
  NOR2_X1 U1177 ( .A1(n180), .A2(n58), .ZN(\ab[14][29] ) );
  NOR2_X1 U1178 ( .A1(n180), .A2(n57), .ZN(\ab[15][29] ) );
  NOR2_X1 U1179 ( .A1(n180), .A2(n56), .ZN(\ab[16][29] ) );
  NOR2_X1 U1180 ( .A1(n180), .A2(n55), .ZN(\ab[17][29] ) );
  AND2_X1 U1181 ( .A1(\SUMB[31][3] ), .A2(\CARRYB[31][2] ), .ZN(\A2[33] ) );
  AND2_X1 U1182 ( .A1(\SUMB[31][5] ), .A2(\CARRYB[31][4] ), .ZN(\A2[35] ) );
  AND2_X1 U1183 ( .A1(\SUMB[31][2] ), .A2(\CARRYB[31][1] ), .ZN(\A2[32] ) );
  AND2_X1 U1184 ( .A1(\SUMB[31][1] ), .A2(\CARRYB[31][0] ), .ZN(\A2[31] ) );
  AND2_X1 U1185 ( .A1(\SUMB[31][7] ), .A2(\CARRYB[31][6] ), .ZN(\A2[37] ) );
  AND2_X1 U1186 ( .A1(\SUMB[31][9] ), .A2(\CARRYB[31][8] ), .ZN(\A2[39] ) );
  AND2_X1 U1187 ( .A1(\SUMB[31][11] ), .A2(\CARRYB[31][10] ), .ZN(\A2[41] ) );
  AND2_X1 U1188 ( .A1(\SUMB[31][13] ), .A2(\CARRYB[31][12] ), .ZN(\A2[43] ) );
  AND2_X1 U1189 ( .A1(\SUMB[31][6] ), .A2(\CARRYB[31][5] ), .ZN(\A2[36] ) );
  AND2_X1 U1190 ( .A1(\SUMB[31][10] ), .A2(\CARRYB[31][9] ), .ZN(\A2[40] ) );
  AND2_X1 U1191 ( .A1(\SUMB[31][14] ), .A2(\CARRYB[31][13] ), .ZN(\A2[44] ) );
  AND2_X1 U1192 ( .A1(n67), .A2(\CARRYB[31][3] ), .ZN(\A2[34] ) );
  AND2_X1 U1193 ( .A1(\SUMB[31][8] ), .A2(\CARRYB[31][7] ), .ZN(\A2[38] ) );
  AND2_X1 U1194 ( .A1(\SUMB[31][12] ), .A2(\CARRYB[31][11] ), .ZN(\A2[42] ) );
  BUF_X1 U1195 ( .A(n2), .Z(n206) );
  BUF_X1 U1196 ( .A(n34), .Z(n120) );
  CLKBUF_X1 U1197 ( .A(n33), .Z(n123) );
  NOR2_X1 U1198 ( .A1(n180), .A2(n40), .ZN(\ab[30][29] ) );
  NOR2_X1 U1199 ( .A1(n180), .A2(n54), .ZN(\ab[18][29] ) );
  NOR2_X1 U1200 ( .A1(n180), .A2(n53), .ZN(\ab[19][29] ) );
  NOR2_X1 U1201 ( .A1(n180), .A2(n51), .ZN(\ab[20][29] ) );
  NOR2_X1 U1202 ( .A1(n180), .A2(n50), .ZN(\ab[21][29] ) );
  NOR2_X1 U1203 ( .A1(n180), .A2(n49), .ZN(\ab[22][29] ) );
  NOR2_X1 U1204 ( .A1(n180), .A2(n48), .ZN(\ab[23][29] ) );
  NOR2_X1 U1205 ( .A1(n180), .A2(n42), .ZN(\ab[29][29] ) );
  NOR2_X1 U1206 ( .A1(n180), .A2(n47), .ZN(\ab[24][29] ) );
  NOR2_X1 U1207 ( .A1(n180), .A2(n46), .ZN(\ab[25][29] ) );
  NOR2_X1 U1208 ( .A1(n180), .A2(n45), .ZN(\ab[26][29] ) );
  NOR2_X1 U1209 ( .A1(n180), .A2(n44), .ZN(\ab[27][29] ) );
  NOR2_X1 U1210 ( .A1(n180), .A2(n43), .ZN(\ab[28][29] ) );
  AND2_X1 U1211 ( .A1(\SUMB[31][20] ), .A2(\CARRYB[31][19] ), .ZN(\A2[50] ) );
  AND2_X1 U1212 ( .A1(\SUMB[31][22] ), .A2(\CARRYB[31][21] ), .ZN(\A2[52] ) );
  AND2_X1 U1213 ( .A1(\SUMB[31][18] ), .A2(\CARRYB[31][17] ), .ZN(\A2[48] ) );
  AND2_X1 U1215 ( .A1(\SUMB[31][30] ), .A2(\CARRYB[31][29] ), .ZN(\A2[60] ) );
  AND2_X1 U1217 ( .A1(\SUMB[31][26] ), .A2(\CARRYB[31][25] ), .ZN(\A2[56] ) );
  AND2_X1 U1218 ( .A1(\SUMB[31][28] ), .A2(\CARRYB[31][27] ), .ZN(\A2[58] ) );
  AND2_X1 U1219 ( .A1(\SUMB[31][15] ), .A2(\CARRYB[31][14] ), .ZN(\A2[45] ) );
  AND2_X1 U1220 ( .A1(\SUMB[31][17] ), .A2(\CARRYB[31][16] ), .ZN(\A2[47] ) );
  AND2_X1 U1221 ( .A1(\SUMB[31][24] ), .A2(\CARRYB[31][23] ), .ZN(\A2[54] ) );
  AND2_X1 U1222 ( .A1(\SUMB[31][21] ), .A2(\CARRYB[31][20] ), .ZN(\A2[51] ) );
  AND2_X1 U1223 ( .A1(\SUMB[31][23] ), .A2(\CARRYB[31][22] ), .ZN(\A2[53] ) );
  AND2_X1 U1224 ( .A1(\SUMB[31][19] ), .A2(\CARRYB[31][18] ), .ZN(\A2[49] ) );
  AND2_X1 U1225 ( .A1(\SUMB[31][29] ), .A2(\CARRYB[31][28] ), .ZN(\A2[59] ) );
  AND2_X1 U1226 ( .A1(\SUMB[31][25] ), .A2(\CARRYB[31][24] ), .ZN(\A2[55] ) );
  AND2_X1 U1227 ( .A1(\SUMB[31][27] ), .A2(\CARRYB[31][26] ), .ZN(\A2[57] ) );
  AND2_X1 U1228 ( .A1(\SUMB[31][16] ), .A2(\CARRYB[31][15] ), .ZN(\A2[46] ) );
  AND2_X1 U1229 ( .A1(\SUMB[31][31] ), .A2(\CARRYB[31][30] ), .ZN(\A2[61] ) );
  BUF_X1 U1230 ( .A(QA), .Z(n210) );
  NOR2_X1 U1231 ( .A1(B[4]), .A2(QA), .ZN(\ab[31][4] ) );
  NOR2_X1 U1232 ( .A1(B[3]), .A2(QA), .ZN(\ab[31][3] ) );
  NOR2_X1 U1233 ( .A1(B[2]), .A2(n210), .ZN(\ab[31][2] ) );
  NOR2_X1 U1234 ( .A1(B[5]), .A2(QA), .ZN(\ab[31][5] ) );
  NOR2_X1 U1235 ( .A1(B[14]), .A2(n210), .ZN(\ab[31][14] ) );
  NOR2_X1 U1236 ( .A1(B[1]), .A2(n210), .ZN(\ab[31][1] ) );
  NOR2_X1 U1237 ( .A1(B[13]), .A2(n210), .ZN(\ab[31][13] ) );
  NOR2_X1 U1238 ( .A1(B[6]), .A2(QA), .ZN(\ab[31][6] ) );
  NOR2_X1 U1239 ( .A1(B[8]), .A2(QA), .ZN(\ab[31][8] ) );
  NOR2_X1 U1240 ( .A1(B[7]), .A2(QA), .ZN(\ab[31][7] ) );
  NOR2_X1 U1241 ( .A1(B[12]), .A2(n210), .ZN(\ab[31][12] ) );
  NOR2_X1 U1242 ( .A1(B[9]), .A2(QA), .ZN(\ab[31][9] ) );
  NOR2_X1 U1243 ( .A1(B[11]), .A2(n210), .ZN(\ab[31][11] ) );
  NOR2_X1 U1244 ( .A1(B[10]), .A2(n210), .ZN(\ab[31][10] ) );
  NOR2_X1 U1245 ( .A1(B[15]), .A2(n210), .ZN(\ab[31][15] ) );
  NOR2_X1 U1246 ( .A1(A[2]), .A2(n209), .ZN(\ab[2][31] ) );
  NOR2_X1 U1247 ( .A1(n185), .A2(n106), .ZN(\ab[3][30] ) );
  NOR2_X1 U1248 ( .A1(A[3]), .A2(n208), .ZN(\ab[3][31] ) );
  NOR2_X1 U1249 ( .A1(n185), .A2(n109), .ZN(\ab[4][30] ) );
  NOR2_X1 U1250 ( .A1(A[4]), .A2(n209), .ZN(\ab[4][31] ) );
  NOR2_X1 U1251 ( .A1(n90), .A2(n111), .ZN(\ab[5][30] ) );
  NOR2_X1 U1252 ( .A1(A[5]), .A2(n208), .ZN(\ab[5][31] ) );
  NOR2_X1 U1253 ( .A1(n185), .A2(n113), .ZN(\ab[6][30] ) );
  NOR2_X1 U1254 ( .A1(A[6]), .A2(n209), .ZN(\ab[6][31] ) );
  NOR2_X1 U1255 ( .A1(n91), .A2(n115), .ZN(\ab[7][30] ) );
  NOR2_X1 U1256 ( .A1(A[7]), .A2(n208), .ZN(\ab[7][31] ) );
  NOR2_X1 U1257 ( .A1(n90), .A2(n118), .ZN(\ab[8][30] ) );
  NOR2_X1 U1258 ( .A1(A[8]), .A2(n209), .ZN(\ab[8][31] ) );
  NOR2_X1 U1259 ( .A1(n206), .A2(n185), .ZN(\ab[9][30] ) );
  NOR2_X1 U1260 ( .A1(A[9]), .A2(n208), .ZN(\ab[9][31] ) );
  NOR2_X1 U1261 ( .A1(n91), .A2(n62), .ZN(\ab[10][30] ) );
  NOR2_X1 U1262 ( .A1(A[10]), .A2(n209), .ZN(\ab[10][31] ) );
  NOR2_X1 U1263 ( .A1(n90), .A2(n61), .ZN(\ab[11][30] ) );
  NOR2_X1 U1264 ( .A1(A[11]), .A2(n208), .ZN(\ab[11][31] ) );
  NOR2_X1 U1265 ( .A1(n185), .A2(n60), .ZN(\ab[12][30] ) );
  NOR2_X1 U1266 ( .A1(A[12]), .A2(n208), .ZN(\ab[12][31] ) );
  NOR2_X1 U1267 ( .A1(n91), .A2(n59), .ZN(\ab[13][30] ) );
  NOR2_X1 U1268 ( .A1(A[13]), .A2(n209), .ZN(\ab[13][31] ) );
  NOR2_X1 U1269 ( .A1(n90), .A2(n58), .ZN(\ab[14][30] ) );
  NOR2_X1 U1270 ( .A1(A[14]), .A2(n208), .ZN(\ab[14][31] ) );
  NOR2_X1 U1271 ( .A1(n91), .A2(n57), .ZN(\ab[15][30] ) );
  NOR2_X1 U1272 ( .A1(A[15]), .A2(n209), .ZN(\ab[15][31] ) );
  NOR2_X1 U1273 ( .A1(n90), .A2(n56), .ZN(\ab[16][30] ) );
  AND2_X1 U1274 ( .A1(\ab[1][30] ), .A2(\ab[0][31] ), .ZN(\CARRYB[1][30] ) );
  NOR2_X1 U1275 ( .A1(B[0]), .A2(n210), .ZN(\ab[31][0] ) );
  INV_X1 U1276 ( .A(B[22]), .ZN(n19) );
  INV_X1 U1277 ( .A(B[21]), .ZN(n20) );
  INV_X1 U1278 ( .A(B[14]), .ZN(n28) );
  INV_X1 U1279 ( .A(B[15]), .ZN(n27) );
  INV_X1 U1280 ( .A(B[23]), .ZN(n18) );
  INV_X1 U1281 ( .A(B[2]), .ZN(n11) );
  INV_X1 U1282 ( .A(B[10]), .ZN(n32) );
  INV_X1 U1283 ( .A(B[13]), .ZN(n29) );
  INV_X1 U1284 ( .A(B[20]), .ZN(n21) );
  INV_X1 U1285 ( .A(B[11]), .ZN(n31) );
  INV_X1 U1286 ( .A(B[12]), .ZN(n30) );
  INV_X1 U1287 ( .A(B[16]), .ZN(n26) );
  INV_X1 U1288 ( .A(B[24]), .ZN(n17) );
  INV_X1 U1289 ( .A(B[19]), .ZN(n23) );
  INV_X1 U1290 ( .A(B[1]), .ZN(n22) );
  INV_X1 U1291 ( .A(B[17]), .ZN(n25) );
  INV_X1 U1292 ( .A(B[18]), .ZN(n24) );
  INV_X1 U1293 ( .A(B[25]), .ZN(n16) );
  INV_X1 U1294 ( .A(B[26]), .ZN(n15) );
  INV_X1 U1295 ( .A(B[27]), .ZN(n14) );
  INV_X1 U1296 ( .A(B[28]), .ZN(n13) );
  INV_X1 U1297 ( .A(B[0]), .ZN(n33) );
  INV_X1 U1298 ( .A(B[29]), .ZN(n12) );
  INV_X1 U1299 ( .A(A[2]), .ZN(n41) );
  INV_X1 U1300 ( .A(A[0]), .ZN(n63) );
  INV_X1 U1301 ( .A(ZB), .ZN(QB) );
  INV_X1 U1302 ( .A(B[5]), .ZN(n7) );
  INV_X1 U1303 ( .A(B[4]), .ZN(n8) );
  INV_X1 U1304 ( .A(B[6]), .ZN(n6) );
  INV_X1 U1305 ( .A(B[7]), .ZN(n5) );
  INV_X1 U1306 ( .A(B[3]), .ZN(n9) );
  INV_X1 U1307 ( .A(B[8]), .ZN(n4) );
  INV_X1 U1308 ( .A(A[3]), .ZN(n39) );
  INV_X1 U1309 ( .A(A[4]), .ZN(n38) );
  INV_X1 U1310 ( .A(A[5]), .ZN(n37) );
  INV_X1 U1311 ( .A(A[6]), .ZN(n36) );
  INV_X1 U1312 ( .A(B[9]), .ZN(n3) );
  NOR2_X1 U1313 ( .A1(A[30]), .A2(n209), .ZN(\ab[30][31] ) );
  NOR2_X1 U1314 ( .A1(n89), .A2(QA), .ZN(\ab[31][30] ) );
  NOR2_X1 U1315 ( .A1(B[21]), .A2(n210), .ZN(\ab[31][21] ) );
  NOR2_X1 U1316 ( .A1(B[20]), .A2(n210), .ZN(\ab[31][20] ) );
  NOR2_X1 U1317 ( .A1(B[22]), .A2(QA), .ZN(\ab[31][22] ) );
  NOR2_X1 U1318 ( .A1(B[19]), .A2(n210), .ZN(\ab[31][19] ) );
  NOR2_X1 U1319 ( .A1(B[23]), .A2(QA), .ZN(\ab[31][23] ) );
  NOR2_X1 U1320 ( .A1(B[18]), .A2(n210), .ZN(\ab[31][18] ) );
  NOR2_X1 U1321 ( .A1(B[24]), .A2(QA), .ZN(\ab[31][24] ) );
  NOR2_X1 U1322 ( .A1(n68), .A2(QA), .ZN(\ab[31][29] ) );
  NOR2_X1 U1323 ( .A1(B[28]), .A2(QA), .ZN(\ab[31][28] ) );
  NOR2_X1 U1324 ( .A1(B[17]), .A2(n210), .ZN(\ab[31][17] ) );
  NOR2_X1 U1325 ( .A1(B[26]), .A2(QA), .ZN(\ab[31][26] ) );
  NOR2_X1 U1326 ( .A1(B[25]), .A2(QA), .ZN(\ab[31][25] ) );
  NOR2_X1 U1327 ( .A1(B[27]), .A2(QA), .ZN(\ab[31][27] ) );
  NOR2_X1 U1328 ( .A1(B[16]), .A2(n210), .ZN(\ab[31][16] ) );
  NOR2_X1 U1329 ( .A1(A[29]), .A2(n208), .ZN(\ab[29][31] ) );
  NOR2_X1 U1330 ( .A1(n185), .A2(n40), .ZN(\ab[30][30] ) );
  NOR2_X1 U1331 ( .A1(A[16]), .A2(n209), .ZN(\ab[16][31] ) );
  NOR2_X1 U1332 ( .A1(n185), .A2(n55), .ZN(\ab[17][30] ) );
  NOR2_X1 U1333 ( .A1(A[20]), .A2(n209), .ZN(\ab[20][31] ) );
  NOR2_X1 U1334 ( .A1(n91), .A2(n50), .ZN(\ab[21][30] ) );
  NOR2_X1 U1335 ( .A1(A[21]), .A2(n208), .ZN(\ab[21][31] ) );
  NOR2_X1 U1336 ( .A1(n90), .A2(n49), .ZN(\ab[22][30] ) );
  NOR2_X1 U1337 ( .A1(A[22]), .A2(n209), .ZN(\ab[22][31] ) );
  NOR2_X1 U1338 ( .A1(n185), .A2(n48), .ZN(\ab[23][30] ) );
  NOR2_X1 U1339 ( .A1(A[23]), .A2(n208), .ZN(\ab[23][31] ) );
  NOR2_X1 U1340 ( .A1(n91), .A2(n47), .ZN(\ab[24][30] ) );
  NOR2_X1 U1341 ( .A1(A[24]), .A2(n209), .ZN(\ab[24][31] ) );
  NOR2_X1 U1342 ( .A1(n90), .A2(n46), .ZN(\ab[25][30] ) );
  NOR2_X1 U1343 ( .A1(A[25]), .A2(n208), .ZN(\ab[25][31] ) );
  NOR2_X1 U1344 ( .A1(n185), .A2(n45), .ZN(\ab[26][30] ) );
  NOR2_X1 U1345 ( .A1(A[28]), .A2(n209), .ZN(\ab[28][31] ) );
  NOR2_X1 U1346 ( .A1(n185), .A2(n42), .ZN(\ab[29][30] ) );
  NOR2_X1 U1347 ( .A1(A[26]), .A2(n209), .ZN(\ab[26][31] ) );
  NOR2_X1 U1348 ( .A1(n91), .A2(n44), .ZN(\ab[27][30] ) );
  NOR2_X1 U1349 ( .A1(A[27]), .A2(n208), .ZN(\ab[27][31] ) );
  NOR2_X1 U1350 ( .A1(n90), .A2(n43), .ZN(\ab[28][30] ) );
  NOR2_X1 U1351 ( .A1(A[17]), .A2(n208), .ZN(\ab[17][31] ) );
  NOR2_X1 U1352 ( .A1(n91), .A2(n54), .ZN(\ab[18][30] ) );
  NOR2_X1 U1353 ( .A1(A[18]), .A2(n209), .ZN(\ab[18][31] ) );
  NOR2_X1 U1354 ( .A1(n90), .A2(n53), .ZN(\ab[19][30] ) );
  NOR2_X1 U1355 ( .A1(A[19]), .A2(n208), .ZN(\ab[19][31] ) );
  NOR2_X1 U1356 ( .A1(n185), .A2(n51), .ZN(\ab[20][30] ) );
  INV_X1 U1357 ( .A(A[7]), .ZN(n35) );
  INV_X1 U1358 ( .A(A[8]), .ZN(n34) );
  INV_X1 U1359 ( .A(A[9]), .ZN(n2) );
  INV_X1 U1360 ( .A(ZA), .ZN(QA) );
  NOR2_X1 U1361 ( .A1(A[1]), .A2(QB), .ZN(\ab[1][31] ) );
  INV_X1 U1362 ( .A(A[1]), .ZN(n52) );
  INV_X1 U1363 ( .A(n66), .ZN(n10) );
endmodule


module Multiplier_NBIT_DATA32_DW02_mult_0 ( A, B, TC, PRODUCT );
  input [31:0] A;
  input [31:0] B;
  output [63:0] PRODUCT;
  input TC;
  wire   \ab[31][30] , \ab[31][29] , \ab[31][28] , \ab[31][27] , \ab[31][26] ,
         \ab[31][25] , \ab[31][24] , \ab[31][23] , \ab[31][22] , \ab[31][21] ,
         \ab[31][20] , \ab[31][19] , \ab[31][18] , \ab[31][17] , \ab[31][16] ,
         \ab[31][15] , \ab[31][14] , \ab[31][13] , \ab[31][12] , \ab[31][11] ,
         \ab[31][10] , \ab[31][9] , \ab[31][8] , \ab[31][7] , \ab[31][6] ,
         \ab[31][5] , \ab[31][4] , \ab[31][3] , \ab[31][2] , \ab[31][1] ,
         \ab[31][0] , \ab[30][31] , \ab[30][30] , \ab[30][29] , \ab[30][28] ,
         \ab[30][27] , \ab[30][26] , \ab[30][25] , \ab[30][24] , \ab[30][23] ,
         \ab[30][22] , \ab[30][21] , \ab[30][20] , \ab[30][19] , \ab[30][18] ,
         \ab[30][17] , \ab[30][16] , \ab[30][15] , \ab[30][14] , \ab[30][13] ,
         \ab[30][12] , \ab[30][11] , \ab[30][10] , \ab[30][9] , \ab[30][8] ,
         \ab[30][7] , \ab[30][6] , \ab[30][5] , \ab[30][4] , \ab[30][3] ,
         \ab[30][2] , \ab[30][1] , \ab[30][0] , \ab[29][31] , \ab[29][30] ,
         \ab[29][29] , \ab[29][28] , \ab[29][27] , \ab[29][26] , \ab[29][25] ,
         \ab[29][24] , \ab[29][23] , \ab[29][22] , \ab[29][21] , \ab[29][20] ,
         \ab[29][19] , \ab[29][18] , \ab[29][17] , \ab[29][16] , \ab[29][15] ,
         \ab[29][14] , \ab[29][13] , \ab[29][12] , \ab[29][11] , \ab[29][10] ,
         \ab[29][9] , \ab[29][8] , \ab[29][7] , \ab[29][6] , \ab[29][5] ,
         \ab[29][4] , \ab[29][3] , \ab[29][2] , \ab[29][1] , \ab[29][0] ,
         \ab[28][31] , \ab[28][30] , \ab[28][29] , \ab[28][28] , \ab[28][27] ,
         \ab[28][26] , \ab[28][25] , \ab[28][24] , \ab[28][23] , \ab[28][22] ,
         \ab[28][21] , \ab[28][20] , \ab[28][19] , \ab[28][18] , \ab[28][17] ,
         \ab[28][16] , \ab[28][15] , \ab[28][14] , \ab[28][13] , \ab[28][12] ,
         \ab[28][11] , \ab[28][10] , \ab[28][9] , \ab[28][8] , \ab[28][7] ,
         \ab[28][6] , \ab[28][5] , \ab[28][4] , \ab[28][3] , \ab[28][2] ,
         \ab[28][1] , \ab[28][0] , \ab[27][31] , \ab[27][30] , \ab[27][29] ,
         \ab[27][28] , \ab[27][27] , \ab[27][26] , \ab[27][25] , \ab[27][24] ,
         \ab[27][23] , \ab[27][22] , \ab[27][21] , \ab[27][20] , \ab[27][19] ,
         \ab[27][18] , \ab[27][17] , \ab[27][16] , \ab[27][15] , \ab[27][14] ,
         \ab[27][13] , \ab[27][12] , \ab[27][11] , \ab[27][10] , \ab[27][9] ,
         \ab[27][8] , \ab[27][7] , \ab[27][6] , \ab[27][5] , \ab[27][4] ,
         \ab[27][3] , \ab[27][2] , \ab[27][1] , \ab[27][0] , \ab[26][31] ,
         \ab[26][30] , \ab[26][29] , \ab[26][28] , \ab[26][27] , \ab[26][26] ,
         \ab[26][25] , \ab[26][24] , \ab[26][23] , \ab[26][22] , \ab[26][21] ,
         \ab[26][20] , \ab[26][19] , \ab[26][18] , \ab[26][17] , \ab[26][16] ,
         \ab[26][15] , \ab[26][14] , \ab[26][13] , \ab[26][12] , \ab[26][11] ,
         \ab[26][10] , \ab[26][9] , \ab[26][8] , \ab[26][7] , \ab[26][6] ,
         \ab[26][5] , \ab[26][4] , \ab[26][3] , \ab[26][2] , \ab[26][1] ,
         \ab[26][0] , \ab[25][31] , \ab[25][30] , \ab[25][29] , \ab[25][28] ,
         \ab[25][27] , \ab[25][26] , \ab[25][25] , \ab[25][24] , \ab[25][23] ,
         \ab[25][22] , \ab[25][21] , \ab[25][20] , \ab[25][19] , \ab[25][18] ,
         \ab[25][17] , \ab[25][16] , \ab[25][15] , \ab[25][14] , \ab[25][13] ,
         \ab[25][12] , \ab[25][11] , \ab[25][10] , \ab[25][9] , \ab[25][8] ,
         \ab[25][7] , \ab[25][6] , \ab[25][5] , \ab[25][4] , \ab[25][3] ,
         \ab[25][2] , \ab[25][1] , \ab[25][0] , \ab[24][31] , \ab[24][30] ,
         \ab[24][29] , \ab[24][28] , \ab[24][27] , \ab[24][26] , \ab[24][25] ,
         \ab[24][24] , \ab[24][23] , \ab[24][22] , \ab[24][21] , \ab[24][20] ,
         \ab[24][19] , \ab[24][18] , \ab[24][17] , \ab[24][16] , \ab[24][15] ,
         \ab[24][14] , \ab[24][13] , \ab[24][12] , \ab[24][11] , \ab[24][10] ,
         \ab[24][9] , \ab[24][8] , \ab[24][7] , \ab[24][6] , \ab[24][5] ,
         \ab[24][4] , \ab[24][3] , \ab[24][2] , \ab[24][1] , \ab[24][0] ,
         \ab[23][31] , \ab[23][30] , \ab[23][29] , \ab[23][28] , \ab[23][27] ,
         \ab[23][26] , \ab[23][25] , \ab[23][24] , \ab[23][23] , \ab[23][22] ,
         \ab[23][21] , \ab[23][20] , \ab[23][19] , \ab[23][18] , \ab[23][17] ,
         \ab[23][16] , \ab[23][15] , \ab[23][14] , \ab[23][13] , \ab[23][12] ,
         \ab[23][11] , \ab[23][10] , \ab[23][9] , \ab[23][8] , \ab[23][7] ,
         \ab[23][6] , \ab[23][5] , \ab[23][4] , \ab[23][3] , \ab[23][2] ,
         \ab[23][1] , \ab[23][0] , \ab[22][31] , \ab[22][30] , \ab[22][29] ,
         \ab[22][28] , \ab[22][27] , \ab[22][26] , \ab[22][25] , \ab[22][24] ,
         \ab[22][23] , \ab[22][22] , \ab[22][21] , \ab[22][20] , \ab[22][19] ,
         \ab[22][18] , \ab[22][17] , \ab[22][16] , \ab[22][15] , \ab[22][14] ,
         \ab[22][13] , \ab[22][12] , \ab[22][11] , \ab[22][10] , \ab[22][9] ,
         \ab[22][8] , \ab[22][7] , \ab[22][6] , \ab[22][5] , \ab[22][4] ,
         \ab[22][3] , \ab[22][2] , \ab[22][1] , \ab[22][0] , \ab[21][31] ,
         \ab[21][30] , \ab[21][29] , \ab[21][28] , \ab[21][27] , \ab[21][26] ,
         \ab[21][25] , \ab[21][24] , \ab[21][23] , \ab[21][22] , \ab[21][21] ,
         \ab[21][20] , \ab[21][19] , \ab[21][18] , \ab[21][17] , \ab[21][16] ,
         \ab[21][15] , \ab[21][14] , \ab[21][13] , \ab[21][12] , \ab[21][11] ,
         \ab[21][10] , \ab[21][9] , \ab[21][8] , \ab[21][7] , \ab[21][6] ,
         \ab[21][5] , \ab[21][4] , \ab[21][3] , \ab[21][2] , \ab[21][1] ,
         \ab[21][0] , \ab[20][31] , \ab[20][30] , \ab[20][29] , \ab[20][28] ,
         \ab[20][27] , \ab[20][26] , \ab[20][25] , \ab[20][24] , \ab[20][23] ,
         \ab[20][22] , \ab[20][21] , \ab[20][20] , \ab[20][19] , \ab[20][18] ,
         \ab[20][17] , \ab[20][16] , \ab[20][15] , \ab[20][14] , \ab[20][13] ,
         \ab[20][12] , \ab[20][11] , \ab[20][10] , \ab[20][9] , \ab[20][8] ,
         \ab[20][7] , \ab[20][6] , \ab[20][5] , \ab[20][4] , \ab[20][3] ,
         \ab[20][2] , \ab[20][1] , \ab[20][0] , \ab[19][31] , \ab[19][30] ,
         \ab[19][29] , \ab[19][28] , \ab[19][27] , \ab[19][26] , \ab[19][25] ,
         \ab[19][24] , \ab[19][23] , \ab[19][22] , \ab[19][21] , \ab[19][20] ,
         \ab[19][19] , \ab[19][18] , \ab[19][17] , \ab[19][16] , \ab[19][15] ,
         \ab[19][14] , \ab[19][13] , \ab[19][12] , \ab[19][11] , \ab[19][10] ,
         \ab[19][9] , \ab[19][8] , \ab[19][7] , \ab[19][6] , \ab[19][5] ,
         \ab[19][4] , \ab[19][3] , \ab[19][2] , \ab[19][1] , \ab[19][0] ,
         \ab[18][31] , \ab[18][30] , \ab[18][29] , \ab[18][28] , \ab[18][27] ,
         \ab[18][26] , \ab[18][25] , \ab[18][24] , \ab[18][23] , \ab[18][22] ,
         \ab[18][21] , \ab[18][20] , \ab[18][19] , \ab[18][18] , \ab[18][17] ,
         \ab[18][16] , \ab[18][15] , \ab[18][14] , \ab[18][13] , \ab[18][12] ,
         \ab[18][11] , \ab[18][10] , \ab[18][9] , \ab[18][8] , \ab[18][7] ,
         \ab[18][6] , \ab[18][5] , \ab[18][4] , \ab[18][3] , \ab[18][2] ,
         \ab[18][1] , \ab[18][0] , \ab[17][31] , \ab[17][30] , \ab[17][29] ,
         \ab[17][28] , \ab[17][27] , \ab[17][26] , \ab[17][25] , \ab[17][24] ,
         \ab[17][23] , \ab[17][22] , \ab[17][21] , \ab[17][20] , \ab[17][19] ,
         \ab[17][18] , \ab[17][17] , \ab[17][16] , \ab[17][15] , \ab[17][14] ,
         \ab[17][13] , \ab[17][12] , \ab[17][11] , \ab[17][10] , \ab[17][9] ,
         \ab[17][8] , \ab[17][7] , \ab[17][6] , \ab[17][5] , \ab[17][4] ,
         \ab[17][3] , \ab[17][2] , \ab[17][1] , \ab[17][0] , \ab[16][31] ,
         \ab[16][30] , \ab[16][29] , \ab[16][28] , \ab[16][27] , \ab[16][26] ,
         \ab[16][25] , \ab[16][24] , \ab[16][23] , \ab[16][22] , \ab[16][21] ,
         \ab[16][20] , \ab[16][19] , \ab[16][18] , \ab[16][17] , \ab[16][16] ,
         \ab[16][15] , \ab[16][14] , \ab[16][13] , \ab[16][12] , \ab[16][11] ,
         \ab[16][10] , \ab[16][9] , \ab[16][8] , \ab[16][7] , \ab[16][6] ,
         \ab[16][5] , \ab[16][4] , \ab[16][3] , \ab[16][2] , \ab[16][1] ,
         \ab[16][0] , \ab[15][31] , \ab[15][30] , \ab[15][29] , \ab[15][28] ,
         \ab[15][27] , \ab[15][26] , \ab[15][25] , \ab[15][24] , \ab[15][23] ,
         \ab[15][22] , \ab[15][21] , \ab[15][20] , \ab[15][19] , \ab[15][18] ,
         \ab[15][17] , \ab[15][16] , \ab[15][15] , \ab[15][14] , \ab[15][13] ,
         \ab[15][12] , \ab[15][11] , \ab[15][10] , \ab[15][9] , \ab[15][8] ,
         \ab[15][7] , \ab[15][6] , \ab[15][5] , \ab[15][4] , \ab[15][3] ,
         \ab[15][2] , \ab[15][1] , \ab[15][0] , \ab[14][31] , \ab[14][30] ,
         \ab[14][29] , \ab[14][28] , \ab[14][27] , \ab[14][26] , \ab[14][25] ,
         \ab[14][24] , \ab[14][23] , \ab[14][22] , \ab[14][21] , \ab[14][20] ,
         \ab[14][19] , \ab[14][18] , \ab[14][17] , \ab[14][16] , \ab[14][15] ,
         \ab[14][14] , \ab[14][13] , \ab[14][12] , \ab[14][11] , \ab[14][10] ,
         \ab[14][9] , \ab[14][8] , \ab[14][7] , \ab[14][6] , \ab[14][5] ,
         \ab[14][4] , \ab[14][3] , \ab[14][2] , \ab[14][1] , \ab[14][0] ,
         \ab[13][31] , \ab[13][30] , \ab[13][29] , \ab[13][28] , \ab[13][27] ,
         \ab[13][26] , \ab[13][25] , \ab[13][24] , \ab[13][23] , \ab[13][22] ,
         \ab[13][21] , \ab[13][20] , \ab[13][19] , \ab[13][18] , \ab[13][17] ,
         \ab[13][16] , \ab[13][15] , \ab[13][14] , \ab[13][13] , \ab[13][12] ,
         \ab[13][11] , \ab[13][10] , \ab[13][9] , \ab[13][8] , \ab[13][7] ,
         \ab[13][6] , \ab[13][5] , \ab[13][4] , \ab[13][3] , \ab[13][2] ,
         \ab[13][1] , \ab[13][0] , \ab[12][31] , \ab[12][30] , \ab[12][29] ,
         \ab[12][28] , \ab[12][27] , \ab[12][26] , \ab[12][25] , \ab[12][24] ,
         \ab[12][23] , \ab[12][22] , \ab[12][21] , \ab[12][20] , \ab[12][19] ,
         \ab[12][18] , \ab[12][17] , \ab[12][16] , \ab[12][15] , \ab[12][14] ,
         \ab[12][13] , \ab[12][12] , \ab[12][11] , \ab[12][10] , \ab[12][9] ,
         \ab[12][8] , \ab[12][7] , \ab[12][6] , \ab[12][5] , \ab[12][4] ,
         \ab[12][3] , \ab[12][2] , \ab[12][1] , \ab[12][0] , \ab[11][31] ,
         \ab[11][30] , \ab[11][29] , \ab[11][28] , \ab[11][27] , \ab[11][26] ,
         \ab[11][25] , \ab[11][24] , \ab[11][23] , \ab[11][22] , \ab[11][21] ,
         \ab[11][20] , \ab[11][19] , \ab[11][18] , \ab[11][17] , \ab[11][16] ,
         \ab[11][15] , \ab[11][14] , \ab[11][13] , \ab[11][12] , \ab[11][11] ,
         \ab[11][10] , \ab[11][9] , \ab[11][8] , \ab[11][7] , \ab[11][6] ,
         \ab[11][5] , \ab[11][4] , \ab[11][3] , \ab[11][2] , \ab[11][1] ,
         \ab[11][0] , \ab[10][31] , \ab[10][30] , \ab[10][29] , \ab[10][28] ,
         \ab[10][27] , \ab[10][26] , \ab[10][25] , \ab[10][24] , \ab[10][23] ,
         \ab[10][22] , \ab[10][21] , \ab[10][20] , \ab[10][19] , \ab[10][18] ,
         \ab[10][17] , \ab[10][16] , \ab[10][15] , \ab[10][14] , \ab[10][13] ,
         \ab[10][12] , \ab[10][11] , \ab[10][10] , \ab[10][9] , \ab[10][8] ,
         \ab[10][7] , \ab[10][6] , \ab[10][5] , \ab[10][4] , \ab[10][3] ,
         \ab[10][2] , \ab[10][1] , \ab[10][0] , \ab[9][31] , \ab[9][30] ,
         \ab[9][29] , \ab[9][28] , \ab[9][27] , \ab[9][26] , \ab[9][25] ,
         \ab[9][24] , \ab[9][23] , \ab[9][22] , \ab[9][21] , \ab[9][20] ,
         \ab[9][19] , \ab[9][18] , \ab[9][17] , \ab[9][16] , \ab[9][15] ,
         \ab[9][14] , \ab[9][13] , \ab[9][12] , \ab[9][11] , \ab[9][10] ,
         \ab[9][9] , \ab[9][8] , \ab[9][7] , \ab[9][6] , \ab[9][5] ,
         \ab[9][4] , \ab[9][3] , \ab[9][2] , \ab[9][1] , \ab[9][0] ,
         \ab[8][31] , \ab[8][30] , \ab[8][29] , \ab[8][28] , \ab[8][27] ,
         \ab[8][26] , \ab[8][25] , \ab[8][24] , \ab[8][23] , \ab[8][22] ,
         \ab[8][21] , \ab[8][20] , \ab[8][19] , \ab[8][18] , \ab[8][17] ,
         \ab[8][16] , \ab[8][15] , \ab[8][14] , \ab[8][13] , \ab[8][12] ,
         \ab[8][11] , \ab[8][10] , \ab[8][9] , \ab[8][8] , \ab[8][7] ,
         \ab[8][6] , \ab[8][5] , \ab[8][4] , \ab[8][3] , \ab[8][2] ,
         \ab[8][1] , \ab[8][0] , \ab[7][31] , \ab[7][30] , \ab[7][29] ,
         \ab[7][28] , \ab[7][27] , \ab[7][26] , \ab[7][25] , \ab[7][24] ,
         \ab[7][23] , \ab[7][22] , \ab[7][21] , \ab[7][20] , \ab[7][19] ,
         \ab[7][18] , \ab[7][17] , \ab[7][16] , \ab[7][15] , \ab[7][14] ,
         \ab[7][13] , \ab[7][12] , \ab[7][11] , \ab[7][10] , \ab[7][9] ,
         \ab[7][8] , \ab[7][7] , \ab[7][6] , \ab[7][5] , \ab[7][4] ,
         \ab[7][3] , \ab[7][2] , \ab[7][1] , \ab[7][0] , \ab[6][31] ,
         \ab[6][30] , \ab[6][29] , \ab[6][28] , \ab[6][27] , \ab[6][26] ,
         \ab[6][25] , \ab[6][24] , \ab[6][23] , \ab[6][22] , \ab[6][21] ,
         \ab[6][20] , \ab[6][19] , \ab[6][18] , \ab[6][17] , \ab[6][16] ,
         \ab[6][15] , \ab[6][14] , \ab[6][13] , \ab[6][12] , \ab[6][11] ,
         \ab[6][10] , \ab[6][9] , \ab[6][8] , \ab[6][7] , \ab[6][6] ,
         \ab[6][5] , \ab[6][4] , \ab[6][3] , \ab[6][2] , \ab[6][1] ,
         \ab[6][0] , \ab[5][31] , \ab[5][30] , \ab[5][29] , \ab[5][28] ,
         \ab[5][27] , \ab[5][26] , \ab[5][25] , \ab[5][24] , \ab[5][23] ,
         \ab[5][22] , \ab[5][21] , \ab[5][20] , \ab[5][19] , \ab[5][18] ,
         \ab[5][17] , \ab[5][16] , \ab[5][15] , \ab[5][14] , \ab[5][13] ,
         \ab[5][12] , \ab[5][11] , \ab[5][10] , \ab[5][9] , \ab[5][8] ,
         \ab[5][7] , \ab[5][6] , \ab[5][5] , \ab[5][4] , \ab[5][3] ,
         \ab[5][2] , \ab[5][1] , \ab[5][0] , \ab[4][31] , \ab[4][30] ,
         \ab[4][29] , \ab[4][28] , \ab[4][27] , \ab[4][26] , \ab[4][25] ,
         \ab[4][24] , \ab[4][23] , \ab[4][22] , \ab[4][21] , \ab[4][20] ,
         \ab[4][19] , \ab[4][18] , \ab[4][17] , \ab[4][16] , \ab[4][15] ,
         \ab[4][14] , \ab[4][13] , \ab[4][12] , \ab[4][11] , \ab[4][10] ,
         \ab[4][9] , \ab[4][8] , \ab[4][7] , \ab[4][6] , \ab[4][5] ,
         \ab[4][4] , \ab[4][3] , \ab[4][2] , \ab[4][1] , \ab[4][0] ,
         \ab[3][31] , \ab[3][30] , \ab[3][29] , \ab[3][28] , \ab[3][27] ,
         \ab[3][26] , \ab[3][25] , \ab[3][24] , \ab[3][23] , \ab[3][22] ,
         \ab[3][21] , \ab[3][20] , \ab[3][19] , \ab[3][18] , \ab[3][17] ,
         \ab[3][16] , \ab[3][15] , \ab[3][14] , \ab[3][13] , \ab[3][12] ,
         \ab[3][11] , \ab[3][10] , \ab[3][9] , \ab[3][8] , \ab[3][7] ,
         \ab[3][6] , \ab[3][5] , \ab[3][4] , \ab[3][3] , \ab[3][2] ,
         \ab[3][1] , \ab[3][0] , \ab[2][31] , \ab[2][29] , \ab[2][28] ,
         \ab[2][27] , \ab[2][26] , \ab[2][25] , \ab[2][24] , \ab[2][23] ,
         \ab[2][22] , \ab[2][21] , \ab[2][20] , \ab[2][19] , \ab[2][18] ,
         \ab[2][17] , \ab[2][16] , \ab[2][15] , \ab[2][14] , \ab[2][13] ,
         \ab[2][12] , \ab[2][11] , \ab[2][10] , \ab[2][9] , \ab[2][8] ,
         \ab[2][7] , \ab[2][6] , \ab[2][5] , \ab[2][4] , \ab[2][3] ,
         \ab[2][2] , \ab[2][1] , \ab[2][0] , \ab[1][29] , \ab[1][28] ,
         \ab[1][27] , \ab[1][26] , \ab[1][25] , \ab[1][24] , \ab[1][23] ,
         \ab[1][22] , \ab[1][21] , \ab[1][20] , \ab[1][19] , \ab[1][18] ,
         \ab[1][17] , \ab[1][16] , \ab[1][15] , \ab[1][14] , \ab[1][13] ,
         \ab[1][12] , \ab[1][11] , \ab[1][10] , \ab[1][9] , \ab[1][8] ,
         \ab[1][7] , \ab[1][6] , \ab[1][5] , \ab[1][4] , \ab[1][3] ,
         \ab[1][2] , \ab[1][1] , \ab[1][0] , \ab[0][30] , \ab[0][29] ,
         \ab[0][28] , \ab[0][27] , \ab[0][26] , \ab[0][25] , \ab[0][24] ,
         \ab[0][23] , \ab[0][22] , \ab[0][21] , \ab[0][20] , \ab[0][19] ,
         \ab[0][18] , \ab[0][17] , \ab[0][16] , \ab[0][15] , \ab[0][14] ,
         \ab[0][13] , \ab[0][12] , \ab[0][11] , \ab[0][10] , \ab[0][9] ,
         \ab[0][8] , \ab[0][7] , \ab[0][6] , \ab[0][5] , \ab[0][4] ,
         \ab[0][3] , \ab[0][2] , \ab[0][1] , \CARRYB[15][30] ,
         \CARRYB[15][29] , \CARRYB[15][28] , \CARRYB[15][27] ,
         \CARRYB[15][26] , \CARRYB[15][25] , \CARRYB[15][24] ,
         \CARRYB[15][23] , \CARRYB[15][22] , \CARRYB[15][21] ,
         \CARRYB[15][20] , \CARRYB[15][16] , \CARRYB[15][15] ,
         \CARRYB[15][14] , \CARRYB[15][13] , \CARRYB[15][12] ,
         \CARRYB[15][11] , \CARRYB[15][10] , \CARRYB[15][9] , \CARRYB[15][8] ,
         \CARRYB[15][7] , \CARRYB[15][6] , \CARRYB[15][5] , \CARRYB[15][4] ,
         \CARRYB[15][3] , \CARRYB[15][2] , \CARRYB[15][1] , \CARRYB[15][0] ,
         \CARRYB[14][30] , \CARRYB[14][29] , \CARRYB[14][28] ,
         \CARRYB[14][27] , \CARRYB[14][26] , \CARRYB[14][25] ,
         \CARRYB[14][24] , \CARRYB[14][23] , \CARRYB[14][22] ,
         \CARRYB[14][21] , \CARRYB[14][17] , \CARRYB[14][16] ,
         \CARRYB[14][15] , \CARRYB[14][14] , \CARRYB[14][13] ,
         \CARRYB[14][12] , \CARRYB[14][11] , \CARRYB[14][10] , \CARRYB[14][9] ,
         \CARRYB[14][8] , \CARRYB[14][7] , \CARRYB[14][6] , \CARRYB[14][5] ,
         \CARRYB[14][4] , \CARRYB[14][3] , \CARRYB[14][2] , \CARRYB[14][1] ,
         \CARRYB[14][0] , \CARRYB[13][30] , \CARRYB[13][29] , \CARRYB[13][28] ,
         \CARRYB[13][27] , \CARRYB[13][26] , \CARRYB[13][25] ,
         \CARRYB[13][24] , \CARRYB[13][23] , \CARRYB[13][22] ,
         \CARRYB[13][18] , \CARRYB[13][17] , \CARRYB[13][16] ,
         \CARRYB[13][15] , \CARRYB[13][14] , \CARRYB[13][13] ,
         \CARRYB[13][12] , \CARRYB[13][11] , \CARRYB[13][10] , \CARRYB[13][9] ,
         \CARRYB[13][8] , \CARRYB[13][7] , \CARRYB[13][6] , \CARRYB[13][5] ,
         \CARRYB[13][4] , \CARRYB[13][3] , \CARRYB[13][2] , \CARRYB[13][1] ,
         \CARRYB[13][0] , \CARRYB[12][30] , \CARRYB[12][29] , \CARRYB[12][28] ,
         \CARRYB[12][27] , \CARRYB[12][26] , \CARRYB[12][25] ,
         \CARRYB[12][24] , \CARRYB[12][23] , \CARRYB[12][19] ,
         \CARRYB[12][18] , \CARRYB[12][17] , \CARRYB[12][16] ,
         \CARRYB[12][15] , \CARRYB[12][14] , \CARRYB[12][13] ,
         \CARRYB[12][12] , \CARRYB[12][11] , \CARRYB[12][10] , \CARRYB[12][9] ,
         \CARRYB[12][8] , \CARRYB[12][7] , \CARRYB[12][6] , \CARRYB[12][5] ,
         \CARRYB[12][4] , \CARRYB[12][3] , \CARRYB[12][2] , \CARRYB[12][1] ,
         \CARRYB[12][0] , \CARRYB[11][30] , \CARRYB[11][29] , \CARRYB[11][28] ,
         \CARRYB[11][27] , \CARRYB[11][26] , \CARRYB[11][25] ,
         \CARRYB[11][24] , \CARRYB[11][20] , \CARRYB[11][19] ,
         \CARRYB[11][18] , \CARRYB[11][17] , \CARRYB[11][16] ,
         \CARRYB[11][15] , \CARRYB[11][14] , \CARRYB[11][13] ,
         \CARRYB[11][12] , \CARRYB[11][11] , \CARRYB[11][10] , \CARRYB[11][9] ,
         \CARRYB[11][8] , \CARRYB[11][7] , \CARRYB[11][6] , \CARRYB[11][5] ,
         \CARRYB[11][4] , \CARRYB[11][3] , \CARRYB[11][2] , \CARRYB[11][1] ,
         \CARRYB[11][0] , \CARRYB[10][30] , \CARRYB[10][29] , \CARRYB[10][28] ,
         \CARRYB[10][27] , \CARRYB[10][26] , \CARRYB[10][25] ,
         \CARRYB[10][21] , \CARRYB[10][20] , \CARRYB[10][19] ,
         \CARRYB[10][18] , \CARRYB[10][17] , \CARRYB[10][16] ,
         \CARRYB[10][15] , \CARRYB[10][14] , \CARRYB[10][13] ,
         \CARRYB[10][12] , \CARRYB[10][11] , \CARRYB[10][10] , \CARRYB[10][9] ,
         \CARRYB[10][8] , \CARRYB[10][7] , \CARRYB[10][6] , \CARRYB[10][5] ,
         \CARRYB[10][4] , \CARRYB[10][3] , \CARRYB[10][2] , \CARRYB[10][1] ,
         \CARRYB[10][0] , \CARRYB[9][30] , \CARRYB[9][29] , \CARRYB[9][28] ,
         \CARRYB[9][27] , \CARRYB[9][26] , \CARRYB[9][22] , \CARRYB[9][21] ,
         \CARRYB[9][20] , \CARRYB[9][19] , \CARRYB[9][18] , \CARRYB[9][17] ,
         \CARRYB[9][16] , \CARRYB[9][15] , \CARRYB[9][14] , \CARRYB[9][13] ,
         \CARRYB[9][12] , \CARRYB[9][11] , \CARRYB[9][10] , \CARRYB[9][9] ,
         \CARRYB[9][8] , \CARRYB[9][7] , \CARRYB[9][6] , \CARRYB[9][5] ,
         \CARRYB[9][4] , \CARRYB[9][3] , \CARRYB[9][2] , \CARRYB[9][1] ,
         \CARRYB[9][0] , \CARRYB[8][30] , \CARRYB[8][29] , \CARRYB[8][28] ,
         \CARRYB[8][27] , \CARRYB[8][23] , \CARRYB[8][22] , \CARRYB[8][21] ,
         \CARRYB[8][20] , \CARRYB[8][19] , \CARRYB[8][18] , \CARRYB[8][17] ,
         \CARRYB[8][16] , \CARRYB[8][15] , \CARRYB[8][14] , \CARRYB[8][13] ,
         \CARRYB[8][12] , \CARRYB[8][11] , \CARRYB[8][10] , \CARRYB[8][9] ,
         \CARRYB[8][8] , \CARRYB[8][7] , \CARRYB[8][6] , \CARRYB[8][5] ,
         \CARRYB[8][4] , \CARRYB[8][3] , \CARRYB[8][2] , \CARRYB[8][1] ,
         \CARRYB[8][0] , \CARRYB[7][30] , \CARRYB[7][29] , \CARRYB[7][28] ,
         \CARRYB[7][24] , \CARRYB[7][23] , \CARRYB[7][22] , \CARRYB[7][21] ,
         \CARRYB[7][20] , \CARRYB[7][19] , \CARRYB[7][18] , \CARRYB[7][17] ,
         \CARRYB[7][16] , \CARRYB[7][15] , \CARRYB[7][14] , \CARRYB[7][13] ,
         \CARRYB[7][12] , \CARRYB[7][11] , \CARRYB[7][10] , \CARRYB[7][9] ,
         \CARRYB[7][8] , \CARRYB[7][7] , \CARRYB[7][6] , \CARRYB[7][5] ,
         \CARRYB[7][4] , \CARRYB[7][3] , \CARRYB[7][2] , \CARRYB[7][1] ,
         \CARRYB[7][0] , \CARRYB[6][30] , \CARRYB[6][29] , \CARRYB[6][25] ,
         \CARRYB[6][24] , \CARRYB[6][23] , \CARRYB[6][22] , \CARRYB[6][21] ,
         \CARRYB[6][20] , \CARRYB[6][19] , \CARRYB[6][18] , \CARRYB[6][17] ,
         \CARRYB[6][16] , \CARRYB[6][15] , \CARRYB[6][14] , \CARRYB[6][13] ,
         \CARRYB[6][12] , \CARRYB[6][11] , \CARRYB[6][10] , \CARRYB[6][9] ,
         \CARRYB[6][8] , \CARRYB[6][7] , \CARRYB[6][6] , \CARRYB[6][5] ,
         \CARRYB[6][4] , \CARRYB[6][3] , \CARRYB[6][2] , \CARRYB[6][1] ,
         \CARRYB[6][0] , \CARRYB[5][30] , \CARRYB[5][29] , \CARRYB[5][26] ,
         \CARRYB[5][25] , \CARRYB[5][24] , \CARRYB[5][23] , \CARRYB[5][22] ,
         \CARRYB[5][21] , \CARRYB[5][20] , \CARRYB[5][19] , \CARRYB[5][18] ,
         \CARRYB[5][17] , \CARRYB[5][16] , \CARRYB[5][15] , \CARRYB[5][14] ,
         \CARRYB[5][13] , \CARRYB[5][12] , \CARRYB[5][11] , \CARRYB[5][10] ,
         \CARRYB[5][9] , \CARRYB[5][8] , \CARRYB[5][7] , \CARRYB[5][6] ,
         \CARRYB[5][5] , \CARRYB[5][4] , \CARRYB[5][3] , \CARRYB[5][2] ,
         \CARRYB[5][1] , \CARRYB[5][0] , \CARRYB[4][30] , \CARRYB[4][29] ,
         \CARRYB[4][27] , \CARRYB[4][26] , \CARRYB[4][25] , \CARRYB[4][24] ,
         \CARRYB[4][23] , \CARRYB[4][22] , \CARRYB[4][21] , \CARRYB[4][20] ,
         \CARRYB[4][19] , \CARRYB[4][18] , \CARRYB[4][17] , \CARRYB[4][16] ,
         \CARRYB[4][15] , \CARRYB[4][14] , \CARRYB[4][13] , \CARRYB[4][12] ,
         \CARRYB[4][11] , \CARRYB[4][10] , \CARRYB[4][9] , \CARRYB[4][8] ,
         \CARRYB[4][7] , \CARRYB[4][6] , \CARRYB[4][5] , \CARRYB[4][4] ,
         \CARRYB[4][3] , \CARRYB[4][2] , \CARRYB[4][1] , \CARRYB[4][0] ,
         \CARRYB[3][30] , \CARRYB[3][28] , \CARRYB[3][27] , \CARRYB[3][26] ,
         \CARRYB[3][25] , \CARRYB[3][24] , \CARRYB[3][23] , \CARRYB[3][22] ,
         \CARRYB[3][21] , \CARRYB[3][20] , \CARRYB[3][19] , \CARRYB[3][18] ,
         \CARRYB[3][17] , \CARRYB[3][16] , \CARRYB[3][15] , \CARRYB[3][14] ,
         \CARRYB[3][13] , \CARRYB[3][12] , \CARRYB[3][11] , \CARRYB[3][10] ,
         \CARRYB[3][9] , \CARRYB[3][8] , \CARRYB[3][7] , \CARRYB[3][6] ,
         \CARRYB[3][5] , \CARRYB[3][4] , \CARRYB[3][3] , \CARRYB[3][2] ,
         \CARRYB[3][1] , \CARRYB[3][0] , \CARRYB[2][29] , \CARRYB[2][28] ,
         \CARRYB[2][27] , \CARRYB[2][26] , \CARRYB[2][25] , \CARRYB[2][24] ,
         \CARRYB[2][23] , \CARRYB[2][22] , \CARRYB[2][21] , \CARRYB[2][20] ,
         \CARRYB[2][19] , \CARRYB[2][18] , \CARRYB[2][17] , \CARRYB[2][16] ,
         \CARRYB[2][15] , \CARRYB[2][14] , \CARRYB[2][13] , \CARRYB[2][12] ,
         \CARRYB[2][11] , \CARRYB[2][10] , \CARRYB[2][9] , \CARRYB[2][8] ,
         \CARRYB[2][7] , \CARRYB[2][6] , \CARRYB[2][5] , \CARRYB[2][4] ,
         \CARRYB[2][3] , \CARRYB[2][2] , \CARRYB[2][1] , \CARRYB[2][0] ,
         \CARRYB[1][29] , \CARRYB[1][28] , \CARRYB[1][27] , \CARRYB[1][26] ,
         \CARRYB[1][25] , \CARRYB[1][24] , \CARRYB[1][23] , \CARRYB[1][22] ,
         \CARRYB[1][21] , \CARRYB[1][20] , \CARRYB[1][19] , \CARRYB[1][18] ,
         \CARRYB[1][17] , \CARRYB[1][16] , \CARRYB[1][15] , \CARRYB[1][14] ,
         \CARRYB[1][13] , \CARRYB[1][12] , \CARRYB[1][11] , \CARRYB[1][10] ,
         \CARRYB[1][9] , \CARRYB[1][8] , \CARRYB[1][7] , \CARRYB[1][6] ,
         \CARRYB[1][5] , \CARRYB[1][4] , \CARRYB[1][3] , \CARRYB[1][2] ,
         \CARRYB[1][1] , \CARRYB[1][0] , \SUMB[15][30] , \SUMB[15][29] ,
         \SUMB[15][28] , \SUMB[15][27] , \SUMB[15][26] , \SUMB[15][25] ,
         \SUMB[15][24] , \SUMB[15][23] , \SUMB[15][22] , \SUMB[15][21] ,
         \SUMB[15][16] , \SUMB[15][15] , \SUMB[15][14] , \SUMB[15][13] ,
         \SUMB[15][12] , \SUMB[15][11] , \SUMB[15][10] , \SUMB[15][9] ,
         \SUMB[15][8] , \SUMB[15][7] , \SUMB[15][6] , \SUMB[15][5] ,
         \SUMB[15][4] , \SUMB[15][3] , \SUMB[15][2] , \SUMB[15][1] ,
         \SUMB[14][30] , \SUMB[14][29] , \SUMB[14][28] , \SUMB[14][27] ,
         \SUMB[14][26] , \SUMB[14][25] , \SUMB[14][24] , \SUMB[14][23] ,
         \SUMB[14][22] , \SUMB[14][17] , \SUMB[14][16] , \SUMB[14][15] ,
         \SUMB[14][14] , \SUMB[14][13] , \SUMB[14][12] , \SUMB[14][11] ,
         \SUMB[14][10] , \SUMB[14][9] , \SUMB[14][8] , \SUMB[14][7] ,
         \SUMB[14][6] , \SUMB[14][5] , \SUMB[14][4] , \SUMB[14][3] ,
         \SUMB[14][2] , \SUMB[14][1] , \SUMB[13][30] , \SUMB[13][29] ,
         \SUMB[13][28] , \SUMB[13][27] , \SUMB[13][26] , \SUMB[13][25] ,
         \SUMB[13][24] , \SUMB[13][23] , \SUMB[13][18] , \SUMB[13][17] ,
         \SUMB[13][16] , \SUMB[13][15] , \SUMB[13][14] , \SUMB[13][13] ,
         \SUMB[13][12] , \SUMB[13][11] , \SUMB[13][10] , \SUMB[13][9] ,
         \SUMB[13][8] , \SUMB[13][7] , \SUMB[13][6] , \SUMB[13][5] ,
         \SUMB[13][4] , \SUMB[13][3] , \SUMB[13][2] , \SUMB[13][1] ,
         \SUMB[12][30] , \SUMB[12][29] , \SUMB[12][28] , \SUMB[12][27] ,
         \SUMB[12][26] , \SUMB[12][25] , \SUMB[12][24] , \SUMB[12][19] ,
         \SUMB[12][18] , \SUMB[12][17] , \SUMB[12][16] , \SUMB[12][15] ,
         \SUMB[12][14] , \SUMB[12][13] , \SUMB[12][12] , \SUMB[12][11] ,
         \SUMB[12][10] , \SUMB[12][9] , \SUMB[12][8] , \SUMB[12][7] ,
         \SUMB[12][6] , \SUMB[12][5] , \SUMB[12][4] , \SUMB[12][3] ,
         \SUMB[12][2] , \SUMB[12][1] , \SUMB[11][30] , \SUMB[11][29] ,
         \SUMB[11][28] , \SUMB[11][27] , \SUMB[11][26] , \SUMB[11][25] ,
         \SUMB[11][20] , \SUMB[11][19] , \SUMB[11][18] , \SUMB[11][17] ,
         \SUMB[11][16] , \SUMB[11][15] , \SUMB[11][14] , \SUMB[11][13] ,
         \SUMB[11][12] , \SUMB[11][11] , \SUMB[11][10] , \SUMB[11][9] ,
         \SUMB[11][8] , \SUMB[11][7] , \SUMB[11][6] , \SUMB[11][5] ,
         \SUMB[11][4] , \SUMB[11][3] , \SUMB[11][2] , \SUMB[11][1] ,
         \SUMB[10][30] , \SUMB[10][29] , \SUMB[10][28] , \SUMB[10][27] ,
         \SUMB[10][26] , \SUMB[10][21] , \SUMB[10][20] , \SUMB[10][19] ,
         \SUMB[10][18] , \SUMB[10][17] , \SUMB[10][16] , \SUMB[10][15] ,
         \SUMB[10][14] , \SUMB[10][13] , \SUMB[10][12] , \SUMB[10][11] ,
         \SUMB[10][10] , \SUMB[10][9] , \SUMB[10][8] , \SUMB[10][7] ,
         \SUMB[10][6] , \SUMB[10][5] , \SUMB[10][4] , \SUMB[10][3] ,
         \SUMB[10][2] , \SUMB[10][1] , \SUMB[9][30] , \SUMB[9][29] ,
         \SUMB[9][28] , \SUMB[9][27] , \SUMB[9][22] , \SUMB[9][21] ,
         \SUMB[9][20] , \SUMB[9][19] , \SUMB[9][18] , \SUMB[9][17] ,
         \SUMB[9][16] , \SUMB[9][15] , \SUMB[9][14] , \SUMB[9][13] ,
         \SUMB[9][12] , \SUMB[9][11] , \SUMB[9][10] , \SUMB[9][9] ,
         \SUMB[9][8] , \SUMB[9][7] , \SUMB[9][6] , \SUMB[9][5] , \SUMB[9][4] ,
         \SUMB[9][3] , \SUMB[9][2] , \SUMB[9][1] , \SUMB[8][30] ,
         \SUMB[8][29] , \SUMB[8][28] , \SUMB[8][23] , \SUMB[8][22] ,
         \SUMB[8][21] , \SUMB[8][20] , \SUMB[8][19] , \SUMB[8][18] ,
         \SUMB[8][17] , \SUMB[8][16] , \SUMB[8][15] , \SUMB[8][14] ,
         \SUMB[8][13] , \SUMB[8][12] , \SUMB[8][11] , \SUMB[8][10] ,
         \SUMB[8][9] , \SUMB[8][8] , \SUMB[8][7] , \SUMB[8][6] , \SUMB[8][5] ,
         \SUMB[8][4] , \SUMB[8][3] , \SUMB[8][2] , \SUMB[8][1] , \SUMB[7][30] ,
         \SUMB[7][29] , \SUMB[7][24] , \SUMB[7][23] , \SUMB[7][22] ,
         \SUMB[7][21] , \SUMB[7][20] , \SUMB[7][19] , \SUMB[7][18] ,
         \SUMB[7][17] , \SUMB[7][16] , \SUMB[7][15] , \SUMB[7][14] ,
         \SUMB[7][13] , \SUMB[7][12] , \SUMB[7][11] , \SUMB[7][10] ,
         \SUMB[7][9] , \SUMB[7][8] , \SUMB[7][7] , \SUMB[7][6] , \SUMB[7][5] ,
         \SUMB[7][4] , \SUMB[7][3] , \SUMB[7][2] , \SUMB[7][1] , \SUMB[6][30] ,
         \SUMB[6][29] , \SUMB[6][25] , \SUMB[6][24] , \SUMB[6][23] ,
         \SUMB[6][22] , \SUMB[6][21] , \SUMB[6][20] , \SUMB[6][19] ,
         \SUMB[6][18] , \SUMB[6][17] , \SUMB[6][16] , \SUMB[6][15] ,
         \SUMB[6][14] , \SUMB[6][13] , \SUMB[6][12] , \SUMB[6][11] ,
         \SUMB[6][10] , \SUMB[6][9] , \SUMB[6][8] , \SUMB[6][7] , \SUMB[6][6] ,
         \SUMB[6][5] , \SUMB[6][4] , \SUMB[6][3] , \SUMB[6][2] , \SUMB[6][1] ,
         \SUMB[5][30] , \SUMB[5][26] , \SUMB[5][25] , \SUMB[5][24] ,
         \SUMB[5][23] , \SUMB[5][22] , \SUMB[5][21] , \SUMB[5][20] ,
         \SUMB[5][19] , \SUMB[5][18] , \SUMB[5][17] , \SUMB[5][16] ,
         \SUMB[5][15] , \SUMB[5][14] , \SUMB[5][13] , \SUMB[5][12] ,
         \SUMB[5][11] , \SUMB[5][10] , \SUMB[5][9] , \SUMB[5][8] ,
         \SUMB[5][7] , \SUMB[5][6] , \SUMB[5][5] , \SUMB[5][4] , \SUMB[5][3] ,
         \SUMB[5][2] , \SUMB[5][1] , \SUMB[4][30] , \SUMB[4][27] ,
         \SUMB[4][26] , \SUMB[4][25] , \SUMB[4][24] , \SUMB[4][23] ,
         \SUMB[4][22] , \SUMB[4][21] , \SUMB[4][20] , \SUMB[4][19] ,
         \SUMB[4][18] , \SUMB[4][17] , \SUMB[4][16] , \SUMB[4][15] ,
         \SUMB[4][14] , \SUMB[4][13] , \SUMB[4][12] , \SUMB[4][11] ,
         \SUMB[4][10] , \SUMB[4][9] , \SUMB[4][8] , \SUMB[4][7] , \SUMB[4][6] ,
         \SUMB[4][5] , \SUMB[4][4] , \SUMB[4][3] , \SUMB[4][2] , \SUMB[4][1] ,
         \SUMB[3][30] , \SUMB[3][28] , \SUMB[3][27] , \SUMB[3][26] ,
         \SUMB[3][25] , \SUMB[3][24] , \SUMB[3][23] , \SUMB[3][22] ,
         \SUMB[3][21] , \SUMB[3][20] , \SUMB[3][19] , \SUMB[3][18] ,
         \SUMB[3][17] , \SUMB[3][16] , \SUMB[3][15] , \SUMB[3][14] ,
         \SUMB[3][13] , \SUMB[3][12] , \SUMB[3][11] , \SUMB[3][10] ,
         \SUMB[3][9] , \SUMB[3][8] , \SUMB[3][7] , \SUMB[3][6] , \SUMB[3][5] ,
         \SUMB[3][4] , \SUMB[3][3] , \SUMB[3][2] , \SUMB[3][1] , \SUMB[2][29] ,
         \SUMB[2][28] , \SUMB[2][27] , \SUMB[2][26] , \SUMB[2][25] ,
         \SUMB[2][24] , \SUMB[2][23] , \SUMB[2][22] , \SUMB[2][21] ,
         \SUMB[2][20] , \SUMB[2][19] , \SUMB[2][18] , \SUMB[2][17] ,
         \SUMB[2][16] , \SUMB[2][15] , \SUMB[2][14] , \SUMB[2][13] ,
         \SUMB[2][12] , \SUMB[2][11] , \SUMB[2][10] , \SUMB[2][9] ,
         \SUMB[2][8] , \SUMB[2][7] , \SUMB[2][6] , \SUMB[2][5] , \SUMB[2][4] ,
         \SUMB[2][3] , \SUMB[2][2] , \SUMB[2][1] , \SUMB[1][30] ,
         \SUMB[1][29] , \SUMB[1][28] , \SUMB[1][27] , \SUMB[1][26] ,
         \SUMB[1][25] , \SUMB[1][24] , \SUMB[1][23] , \SUMB[1][22] ,
         \SUMB[1][21] , \SUMB[1][20] , \SUMB[1][19] , \SUMB[1][18] ,
         \SUMB[1][17] , \SUMB[1][16] , \SUMB[1][15] , \SUMB[1][14] ,
         \SUMB[1][13] , \SUMB[1][12] , \SUMB[1][11] , \SUMB[1][10] ,
         \SUMB[1][9] , \SUMB[1][8] , \SUMB[1][7] , \SUMB[1][6] , \SUMB[1][5] ,
         \SUMB[1][4] , \SUMB[1][3] , \SUMB[1][2] , \SUMB[1][1] ,
         \CARRYB[31][30] , \CARRYB[31][29] , \CARRYB[31][28] ,
         \CARRYB[31][27] , \CARRYB[31][26] , \CARRYB[31][25] ,
         \CARRYB[31][24] , \CARRYB[31][23] , \CARRYB[31][22] ,
         \CARRYB[31][21] , \CARRYB[31][20] , \CARRYB[31][19] ,
         \CARRYB[31][18] , \CARRYB[31][17] , \CARRYB[31][16] ,
         \CARRYB[31][15] , \CARRYB[31][14] , \CARRYB[31][13] ,
         \CARRYB[31][12] , \CARRYB[31][11] , \CARRYB[31][10] , \CARRYB[31][9] ,
         \CARRYB[31][8] , \CARRYB[31][7] , \CARRYB[31][6] , \CARRYB[31][5] ,
         \CARRYB[31][4] , \CARRYB[31][2] , \CARRYB[31][1] , \CARRYB[31][0] ,
         \CARRYB[30][30] , \CARRYB[30][29] , \CARRYB[30][28] ,
         \CARRYB[30][27] , \CARRYB[30][26] , \CARRYB[30][25] ,
         \CARRYB[30][24] , \CARRYB[30][23] , \CARRYB[30][22] ,
         \CARRYB[30][21] , \CARRYB[30][20] , \CARRYB[30][19] ,
         \CARRYB[30][18] , \CARRYB[30][17] , \CARRYB[30][16] ,
         \CARRYB[30][15] , \CARRYB[30][14] , \CARRYB[30][13] ,
         \CARRYB[30][12] , \CARRYB[30][11] , \CARRYB[30][10] , \CARRYB[30][9] ,
         \CARRYB[30][8] , \CARRYB[30][7] , \CARRYB[30][6] , \CARRYB[30][5] ,
         \CARRYB[30][3] , \CARRYB[30][2] , \CARRYB[30][1] , \CARRYB[30][0] ,
         \CARRYB[29][30] , \CARRYB[29][29] , \CARRYB[29][28] ,
         \CARRYB[29][27] , \CARRYB[29][26] , \CARRYB[29][25] ,
         \CARRYB[29][24] , \CARRYB[29][23] , \CARRYB[29][22] ,
         \CARRYB[29][21] , \CARRYB[29][20] , \CARRYB[29][19] ,
         \CARRYB[29][18] , \CARRYB[29][17] , \CARRYB[29][16] ,
         \CARRYB[29][15] , \CARRYB[29][14] , \CARRYB[29][13] ,
         \CARRYB[29][12] , \CARRYB[29][11] , \CARRYB[29][10] , \CARRYB[29][9] ,
         \CARRYB[29][8] , \CARRYB[29][7] , \CARRYB[29][6] , \CARRYB[29][4] ,
         \CARRYB[29][3] , \CARRYB[29][2] , \CARRYB[29][1] , \CARRYB[29][0] ,
         \CARRYB[28][30] , \CARRYB[28][29] , \CARRYB[28][28] ,
         \CARRYB[28][27] , \CARRYB[28][26] , \CARRYB[28][25] ,
         \CARRYB[28][24] , \CARRYB[28][23] , \CARRYB[28][22] ,
         \CARRYB[28][21] , \CARRYB[28][20] , \CARRYB[28][19] ,
         \CARRYB[28][18] , \CARRYB[28][17] , \CARRYB[28][16] ,
         \CARRYB[28][15] , \CARRYB[28][14] , \CARRYB[28][13] ,
         \CARRYB[28][12] , \CARRYB[28][11] , \CARRYB[28][10] , \CARRYB[28][9] ,
         \CARRYB[28][8] , \CARRYB[28][7] , \CARRYB[28][5] , \CARRYB[28][4] ,
         \CARRYB[28][3] , \CARRYB[28][2] , \CARRYB[28][1] , \CARRYB[28][0] ,
         \CARRYB[27][30] , \CARRYB[27][29] , \CARRYB[27][28] ,
         \CARRYB[27][27] , \CARRYB[27][26] , \CARRYB[27][25] ,
         \CARRYB[27][24] , \CARRYB[27][23] , \CARRYB[27][22] ,
         \CARRYB[27][21] , \CARRYB[27][20] , \CARRYB[27][19] ,
         \CARRYB[27][18] , \CARRYB[27][17] , \CARRYB[27][16] ,
         \CARRYB[27][15] , \CARRYB[27][14] , \CARRYB[27][13] ,
         \CARRYB[27][12] , \CARRYB[27][11] , \CARRYB[27][10] , \CARRYB[27][9] ,
         \CARRYB[27][8] , \CARRYB[27][6] , \CARRYB[27][5] , \CARRYB[27][4] ,
         \CARRYB[27][3] , \CARRYB[27][2] , \CARRYB[27][1] , \CARRYB[27][0] ,
         \CARRYB[26][30] , \CARRYB[26][29] , \CARRYB[26][28] ,
         \CARRYB[26][27] , \CARRYB[26][26] , \CARRYB[26][25] ,
         \CARRYB[26][24] , \CARRYB[26][23] , \CARRYB[26][22] ,
         \CARRYB[26][21] , \CARRYB[26][20] , \CARRYB[26][19] ,
         \CARRYB[26][18] , \CARRYB[26][17] , \CARRYB[26][16] ,
         \CARRYB[26][15] , \CARRYB[26][14] , \CARRYB[26][13] ,
         \CARRYB[26][12] , \CARRYB[26][11] , \CARRYB[26][10] , \CARRYB[26][9] ,
         \CARRYB[26][7] , \CARRYB[26][6] , \CARRYB[26][5] , \CARRYB[26][4] ,
         \CARRYB[26][3] , \CARRYB[26][2] , \CARRYB[26][1] , \CARRYB[26][0] ,
         \CARRYB[25][30] , \CARRYB[25][29] , \CARRYB[25][28] ,
         \CARRYB[25][27] , \CARRYB[25][26] , \CARRYB[25][25] ,
         \CARRYB[25][24] , \CARRYB[25][23] , \CARRYB[25][22] ,
         \CARRYB[25][21] , \CARRYB[25][20] , \CARRYB[25][19] ,
         \CARRYB[25][18] , \CARRYB[25][17] , \CARRYB[25][16] ,
         \CARRYB[25][15] , \CARRYB[25][14] , \CARRYB[25][13] ,
         \CARRYB[25][12] , \CARRYB[25][11] , \CARRYB[25][10] , \CARRYB[25][8] ,
         \CARRYB[25][7] , \CARRYB[25][6] , \CARRYB[25][5] , \CARRYB[25][4] ,
         \CARRYB[25][3] , \CARRYB[25][2] , \CARRYB[25][1] , \CARRYB[25][0] ,
         \CARRYB[24][30] , \CARRYB[24][29] , \CARRYB[24][28] ,
         \CARRYB[24][27] , \CARRYB[24][26] , \CARRYB[24][25] ,
         \CARRYB[24][24] , \CARRYB[24][23] , \CARRYB[24][22] ,
         \CARRYB[24][21] , \CARRYB[24][20] , \CARRYB[24][19] ,
         \CARRYB[24][18] , \CARRYB[24][17] , \CARRYB[24][16] ,
         \CARRYB[24][15] , \CARRYB[24][14] , \CARRYB[24][13] ,
         \CARRYB[24][12] , \CARRYB[24][11] , \CARRYB[24][9] , \CARRYB[24][8] ,
         \CARRYB[24][7] , \CARRYB[24][6] , \CARRYB[24][5] , \CARRYB[24][4] ,
         \CARRYB[24][3] , \CARRYB[24][2] , \CARRYB[24][1] , \CARRYB[24][0] ,
         \CARRYB[23][30] , \CARRYB[23][29] , \CARRYB[23][28] ,
         \CARRYB[23][27] , \CARRYB[23][26] , \CARRYB[23][25] ,
         \CARRYB[23][24] , \CARRYB[23][23] , \CARRYB[23][22] ,
         \CARRYB[23][21] , \CARRYB[23][20] , \CARRYB[23][19] ,
         \CARRYB[23][18] , \CARRYB[23][17] , \CARRYB[23][16] ,
         \CARRYB[23][15] , \CARRYB[23][14] , \CARRYB[23][13] ,
         \CARRYB[23][12] , \CARRYB[23][10] , \CARRYB[23][9] , \CARRYB[23][8] ,
         \CARRYB[23][7] , \CARRYB[23][6] , \CARRYB[23][5] , \CARRYB[23][4] ,
         \CARRYB[23][3] , \CARRYB[23][2] , \CARRYB[23][1] , \CARRYB[23][0] ,
         \CARRYB[22][30] , \CARRYB[22][29] , \CARRYB[22][28] ,
         \CARRYB[22][27] , \CARRYB[22][26] , \CARRYB[22][25] ,
         \CARRYB[22][24] , \CARRYB[22][23] , \CARRYB[22][22] ,
         \CARRYB[22][21] , \CARRYB[22][20] , \CARRYB[22][19] ,
         \CARRYB[22][18] , \CARRYB[22][17] , \CARRYB[22][16] ,
         \CARRYB[22][15] , \CARRYB[22][14] , \CARRYB[22][13] ,
         \CARRYB[22][11] , \CARRYB[22][10] , \CARRYB[22][9] , \CARRYB[22][8] ,
         \CARRYB[22][7] , \CARRYB[22][6] , \CARRYB[22][5] , \CARRYB[22][4] ,
         \CARRYB[22][3] , \CARRYB[22][2] , \CARRYB[22][1] , \CARRYB[22][0] ,
         \CARRYB[21][30] , \CARRYB[21][29] , \CARRYB[21][28] ,
         \CARRYB[21][27] , \CARRYB[21][26] , \CARRYB[21][25] ,
         \CARRYB[21][24] , \CARRYB[21][23] , \CARRYB[21][22] ,
         \CARRYB[21][21] , \CARRYB[21][20] , \CARRYB[21][19] ,
         \CARRYB[21][18] , \CARRYB[21][17] , \CARRYB[21][16] ,
         \CARRYB[21][15] , \CARRYB[21][14] , \CARRYB[21][12] ,
         \CARRYB[21][11] , \CARRYB[21][10] , \CARRYB[21][9] , \CARRYB[21][8] ,
         \CARRYB[21][7] , \CARRYB[21][6] , \CARRYB[21][5] , \CARRYB[21][4] ,
         \CARRYB[21][3] , \CARRYB[21][2] , \CARRYB[21][1] , \CARRYB[21][0] ,
         \CARRYB[20][30] , \CARRYB[20][29] , \CARRYB[20][28] ,
         \CARRYB[20][27] , \CARRYB[20][26] , \CARRYB[20][25] ,
         \CARRYB[20][24] , \CARRYB[20][23] , \CARRYB[20][22] ,
         \CARRYB[20][21] , \CARRYB[20][20] , \CARRYB[20][19] ,
         \CARRYB[20][18] , \CARRYB[20][17] , \CARRYB[20][16] ,
         \CARRYB[20][15] , \CARRYB[20][13] , \CARRYB[20][12] ,
         \CARRYB[20][11] , \CARRYB[20][10] , \CARRYB[20][9] , \CARRYB[20][8] ,
         \CARRYB[20][7] , \CARRYB[20][6] , \CARRYB[20][5] , \CARRYB[20][4] ,
         \CARRYB[20][3] , \CARRYB[20][2] , \CARRYB[20][1] , \CARRYB[20][0] ,
         \CARRYB[19][30] , \CARRYB[19][29] , \CARRYB[19][28] ,
         \CARRYB[19][27] , \CARRYB[19][26] , \CARRYB[19][25] ,
         \CARRYB[19][24] , \CARRYB[19][23] , \CARRYB[19][22] ,
         \CARRYB[19][21] , \CARRYB[19][20] , \CARRYB[19][19] ,
         \CARRYB[19][18] , \CARRYB[19][17] , \CARRYB[19][16] ,
         \CARRYB[19][14] , \CARRYB[19][13] , \CARRYB[19][12] ,
         \CARRYB[19][11] , \CARRYB[19][10] , \CARRYB[19][9] , \CARRYB[19][8] ,
         \CARRYB[19][7] , \CARRYB[19][6] , \CARRYB[19][5] , \CARRYB[19][4] ,
         \CARRYB[19][3] , \CARRYB[19][2] , \CARRYB[19][1] , \CARRYB[19][0] ,
         \CARRYB[18][30] , \CARRYB[18][29] , \CARRYB[18][28] ,
         \CARRYB[18][27] , \CARRYB[18][26] , \CARRYB[18][25] ,
         \CARRYB[18][24] , \CARRYB[18][23] , \CARRYB[18][22] ,
         \CARRYB[18][21] , \CARRYB[18][20] , \CARRYB[18][19] ,
         \CARRYB[18][18] , \CARRYB[18][17] , \CARRYB[18][14] ,
         \CARRYB[18][13] , \CARRYB[18][12] , \CARRYB[18][11] ,
         \CARRYB[18][10] , \CARRYB[18][9] , \CARRYB[18][8] , \CARRYB[18][7] ,
         \CARRYB[18][6] , \CARRYB[18][5] , \CARRYB[18][4] , \CARRYB[18][3] ,
         \CARRYB[18][2] , \CARRYB[18][1] , \CARRYB[18][0] , \CARRYB[17][30] ,
         \CARRYB[17][29] , \CARRYB[17][28] , \CARRYB[17][27] ,
         \CARRYB[17][26] , \CARRYB[17][25] , \CARRYB[17][24] ,
         \CARRYB[17][23] , \CARRYB[17][22] , \CARRYB[17][21] ,
         \CARRYB[17][20] , \CARRYB[17][19] , \CARRYB[17][18] ,
         \CARRYB[17][14] , \CARRYB[17][13] , \CARRYB[17][12] ,
         \CARRYB[17][11] , \CARRYB[17][10] , \CARRYB[17][9] , \CARRYB[17][8] ,
         \CARRYB[17][7] , \CARRYB[17][6] , \CARRYB[17][5] , \CARRYB[17][4] ,
         \CARRYB[17][3] , \CARRYB[17][2] , \CARRYB[17][1] , \CARRYB[17][0] ,
         \CARRYB[16][30] , \CARRYB[16][29] , \CARRYB[16][28] ,
         \CARRYB[16][27] , \CARRYB[16][26] , \CARRYB[16][25] ,
         \CARRYB[16][24] , \CARRYB[16][23] , \CARRYB[16][22] ,
         \CARRYB[16][21] , \CARRYB[16][20] , \CARRYB[16][19] ,
         \CARRYB[16][15] , \CARRYB[16][14] , \CARRYB[16][13] ,
         \CARRYB[16][12] , \CARRYB[16][11] , \CARRYB[16][10] , \CARRYB[16][9] ,
         \CARRYB[16][8] , \CARRYB[16][7] , \CARRYB[16][6] , \CARRYB[16][5] ,
         \CARRYB[16][4] , \CARRYB[16][3] , \CARRYB[16][2] , \CARRYB[16][1] ,
         \CARRYB[16][0] , \SUMB[31][31] , \SUMB[31][30] , \SUMB[31][29] ,
         \SUMB[31][28] , \SUMB[31][27] , \SUMB[31][26] , \SUMB[31][25] ,
         \SUMB[31][24] , \SUMB[31][23] , \SUMB[31][22] , \SUMB[31][21] ,
         \SUMB[31][20] , \SUMB[31][19] , \SUMB[31][18] , \SUMB[31][17] ,
         \SUMB[31][16] , \SUMB[31][15] , \SUMB[31][14] , \SUMB[31][13] ,
         \SUMB[31][12] , \SUMB[31][11] , \SUMB[31][10] , \SUMB[31][9] ,
         \SUMB[31][8] , \SUMB[31][7] , \SUMB[31][6] , \SUMB[31][5] ,
         \SUMB[31][2] , \SUMB[31][1] , \SUMB[30][30] , \SUMB[30][29] ,
         \SUMB[30][28] , \SUMB[30][27] , \SUMB[30][26] , \SUMB[30][25] ,
         \SUMB[30][24] , \SUMB[30][23] , \SUMB[30][22] , \SUMB[30][21] ,
         \SUMB[30][20] , \SUMB[30][19] , \SUMB[30][18] , \SUMB[30][17] ,
         \SUMB[30][16] , \SUMB[30][15] , \SUMB[30][14] , \SUMB[30][13] ,
         \SUMB[30][12] , \SUMB[30][11] , \SUMB[30][10] , \SUMB[30][9] ,
         \SUMB[30][8] , \SUMB[30][7] , \SUMB[30][6] , \SUMB[30][3] ,
         \SUMB[30][2] , \SUMB[30][1] , \SUMB[29][30] , \SUMB[29][29] ,
         \SUMB[29][28] , \SUMB[29][27] , \SUMB[29][26] , \SUMB[29][25] ,
         \SUMB[29][24] , \SUMB[29][23] , \SUMB[29][22] , \SUMB[29][21] ,
         \SUMB[29][20] , \SUMB[29][19] , \SUMB[29][18] , \SUMB[29][17] ,
         \SUMB[29][16] , \SUMB[29][15] , \SUMB[29][14] , \SUMB[29][13] ,
         \SUMB[29][12] , \SUMB[29][11] , \SUMB[29][10] , \SUMB[29][9] ,
         \SUMB[29][8] , \SUMB[29][7] , \SUMB[29][4] , \SUMB[29][3] ,
         \SUMB[29][2] , \SUMB[29][1] , \SUMB[28][30] , \SUMB[28][29] ,
         \SUMB[28][28] , \SUMB[28][27] , \SUMB[28][26] , \SUMB[28][25] ,
         \SUMB[28][24] , \SUMB[28][23] , \SUMB[28][22] , \SUMB[28][21] ,
         \SUMB[28][20] , \SUMB[28][19] , \SUMB[28][18] , \SUMB[28][17] ,
         \SUMB[28][16] , \SUMB[28][15] , \SUMB[28][14] , \SUMB[28][13] ,
         \SUMB[28][12] , \SUMB[28][11] , \SUMB[28][10] , \SUMB[28][9] ,
         \SUMB[28][8] , \SUMB[28][5] , \SUMB[28][4] , \SUMB[28][3] ,
         \SUMB[28][2] , \SUMB[28][1] , \SUMB[27][30] , \SUMB[27][29] ,
         \SUMB[27][28] , \SUMB[27][27] , \SUMB[27][26] , \SUMB[27][25] ,
         \SUMB[27][24] , \SUMB[27][23] , \SUMB[27][22] , \SUMB[27][21] ,
         \SUMB[27][20] , \SUMB[27][19] , \SUMB[27][18] , \SUMB[27][17] ,
         \SUMB[27][16] , \SUMB[27][15] , \SUMB[27][14] , \SUMB[27][13] ,
         \SUMB[27][12] , \SUMB[27][11] , \SUMB[27][10] , \SUMB[27][9] ,
         \SUMB[27][6] , \SUMB[27][5] , \SUMB[27][4] , \SUMB[27][3] ,
         \SUMB[27][2] , \SUMB[27][1] , \SUMB[26][30] , \SUMB[26][29] ,
         \SUMB[26][28] , \SUMB[26][27] , \SUMB[26][26] , \SUMB[26][25] ,
         \SUMB[26][24] , \SUMB[26][23] , \SUMB[26][22] , \SUMB[26][21] ,
         \SUMB[26][20] , \SUMB[26][19] , \SUMB[26][18] , \SUMB[26][17] ,
         \SUMB[26][16] , \SUMB[26][15] , \SUMB[26][14] , \SUMB[26][13] ,
         \SUMB[26][12] , \SUMB[26][11] , \SUMB[26][10] , \SUMB[26][7] ,
         \SUMB[26][6] , \SUMB[26][5] , \SUMB[26][4] , \SUMB[26][3] ,
         \SUMB[26][2] , \SUMB[26][1] , \SUMB[25][30] , \SUMB[25][29] ,
         \SUMB[25][28] , \SUMB[25][27] , \SUMB[25][26] , \SUMB[25][25] ,
         \SUMB[25][24] , \SUMB[25][23] , \SUMB[25][22] , \SUMB[25][21] ,
         \SUMB[25][20] , \SUMB[25][19] , \SUMB[25][18] , \SUMB[25][17] ,
         \SUMB[25][16] , \SUMB[25][15] , \SUMB[25][14] , \SUMB[25][13] ,
         \SUMB[25][12] , \SUMB[25][11] , \SUMB[25][8] , \SUMB[25][7] ,
         \SUMB[25][6] , \SUMB[25][5] , \SUMB[25][4] , \SUMB[25][3] ,
         \SUMB[25][2] , \SUMB[25][1] , \SUMB[24][30] , \SUMB[24][29] ,
         \SUMB[24][28] , \SUMB[24][27] , \SUMB[24][26] , \SUMB[24][25] ,
         \SUMB[24][24] , \SUMB[24][23] , \SUMB[24][22] , \SUMB[24][21] ,
         \SUMB[24][20] , \SUMB[24][19] , \SUMB[24][18] , \SUMB[24][17] ,
         \SUMB[24][16] , \SUMB[24][15] , \SUMB[24][14] , \SUMB[24][13] ,
         \SUMB[24][12] , \SUMB[24][9] , \SUMB[24][8] , \SUMB[24][7] ,
         \SUMB[24][6] , \SUMB[24][5] , \SUMB[24][4] , \SUMB[24][3] ,
         \SUMB[24][2] , \SUMB[24][1] , \SUMB[23][30] , \SUMB[23][29] ,
         \SUMB[23][28] , \SUMB[23][27] , \SUMB[23][26] , \SUMB[23][25] ,
         \SUMB[23][24] , \SUMB[23][23] , \SUMB[23][22] , \SUMB[23][21] ,
         \SUMB[23][20] , \SUMB[23][19] , \SUMB[23][18] , \SUMB[23][17] ,
         \SUMB[23][16] , \SUMB[23][15] , \SUMB[23][14] , \SUMB[23][13] ,
         \SUMB[23][10] , \SUMB[23][9] , \SUMB[23][8] , \SUMB[23][7] ,
         \SUMB[23][6] , \SUMB[23][5] , \SUMB[23][4] , \SUMB[23][3] ,
         \SUMB[23][2] , \SUMB[23][1] , \SUMB[22][30] , \SUMB[22][29] ,
         \SUMB[22][28] , \SUMB[22][27] , \SUMB[22][26] , \SUMB[22][25] ,
         \SUMB[22][24] , \SUMB[22][23] , \SUMB[22][22] , \SUMB[22][21] ,
         \SUMB[22][20] , \SUMB[22][19] , \SUMB[22][18] , \SUMB[22][17] ,
         \SUMB[22][16] , \SUMB[22][15] , \SUMB[22][14] , \SUMB[22][11] ,
         \SUMB[22][10] , \SUMB[22][9] , \SUMB[22][8] , \SUMB[22][7] ,
         \SUMB[22][6] , \SUMB[22][5] , \SUMB[22][4] , \SUMB[22][3] ,
         \SUMB[22][2] , \SUMB[22][1] , \SUMB[21][30] , \SUMB[21][29] ,
         \SUMB[21][28] , \SUMB[21][27] , \SUMB[21][26] , \SUMB[21][25] ,
         \SUMB[21][24] , \SUMB[21][23] , \SUMB[21][22] , \SUMB[21][21] ,
         \SUMB[21][20] , \SUMB[21][19] , \SUMB[21][18] , \SUMB[21][17] ,
         \SUMB[21][16] , \SUMB[21][15] , \SUMB[21][12] , \SUMB[21][11] ,
         \SUMB[21][10] , \SUMB[21][9] , \SUMB[21][8] , \SUMB[21][7] ,
         \SUMB[21][6] , \SUMB[21][5] , \SUMB[21][4] , \SUMB[21][3] ,
         \SUMB[21][2] , \SUMB[21][1] , \SUMB[20][30] , \SUMB[20][29] ,
         \SUMB[20][28] , \SUMB[20][27] , \SUMB[20][26] , \SUMB[20][25] ,
         \SUMB[20][24] , \SUMB[20][23] , \SUMB[20][22] , \SUMB[20][21] ,
         \SUMB[20][20] , \SUMB[20][19] , \SUMB[20][18] , \SUMB[20][17] ,
         \SUMB[20][16] , \SUMB[20][13] , \SUMB[20][12] , \SUMB[20][11] ,
         \SUMB[20][10] , \SUMB[20][9] , \SUMB[20][8] , \SUMB[20][7] ,
         \SUMB[20][6] , \SUMB[20][5] , \SUMB[20][4] , \SUMB[20][3] ,
         \SUMB[20][2] , \SUMB[20][1] , \SUMB[19][30] , \SUMB[19][29] ,
         \SUMB[19][28] , \SUMB[19][27] , \SUMB[19][26] , \SUMB[19][25] ,
         \SUMB[19][24] , \SUMB[19][23] , \SUMB[19][22] , \SUMB[19][21] ,
         \SUMB[19][20] , \SUMB[19][19] , \SUMB[19][18] , \SUMB[19][17] ,
         \SUMB[19][14] , \SUMB[19][13] , \SUMB[19][12] , \SUMB[19][11] ,
         \SUMB[19][10] , \SUMB[19][9] , \SUMB[19][8] , \SUMB[19][7] ,
         \SUMB[19][6] , \SUMB[19][5] , \SUMB[19][4] , \SUMB[19][3] ,
         \SUMB[19][2] , \SUMB[19][1] , \SUMB[18][30] , \SUMB[18][29] ,
         \SUMB[18][28] , \SUMB[18][27] , \SUMB[18][26] , \SUMB[18][25] ,
         \SUMB[18][24] , \SUMB[18][23] , \SUMB[18][22] , \SUMB[18][21] ,
         \SUMB[18][20] , \SUMB[18][19] , \SUMB[18][18] , \SUMB[18][14] ,
         \SUMB[18][13] , \SUMB[18][12] , \SUMB[18][11] , \SUMB[18][10] ,
         \SUMB[18][9] , \SUMB[18][8] , \SUMB[18][7] , \SUMB[18][6] ,
         \SUMB[18][5] , \SUMB[18][4] , \SUMB[18][3] , \SUMB[18][2] ,
         \SUMB[18][1] , \SUMB[17][30] , \SUMB[17][29] , \SUMB[17][28] ,
         \SUMB[17][27] , \SUMB[17][26] , \SUMB[17][25] , \SUMB[17][24] ,
         \SUMB[17][23] , \SUMB[17][22] , \SUMB[17][21] , \SUMB[17][20] ,
         \SUMB[17][19] , \SUMB[17][14] , \SUMB[17][13] , \SUMB[17][12] ,
         \SUMB[17][11] , \SUMB[17][10] , \SUMB[17][9] , \SUMB[17][8] ,
         \SUMB[17][7] , \SUMB[17][6] , \SUMB[17][5] , \SUMB[17][4] ,
         \SUMB[17][3] , \SUMB[17][2] , \SUMB[17][1] , \SUMB[16][30] ,
         \SUMB[16][29] , \SUMB[16][28] , \SUMB[16][27] , \SUMB[16][26] ,
         \SUMB[16][25] , \SUMB[16][24] , \SUMB[16][23] , \SUMB[16][22] ,
         \SUMB[16][21] , \SUMB[16][20] , \SUMB[16][15] , \SUMB[16][14] ,
         \SUMB[16][13] , \SUMB[16][12] , \SUMB[16][11] , \SUMB[16][10] ,
         \SUMB[16][9] , \SUMB[16][8] , \SUMB[16][7] , \SUMB[16][6] ,
         \SUMB[16][5] , \SUMB[16][4] , \SUMB[16][3] , \SUMB[16][2] ,
         \SUMB[16][1] , \A1[60] , \A1[59] , \A1[58] , \A1[57] , \A1[56] ,
         \A1[55] , \A1[54] , \A1[53] , \A1[52] , \A1[51] , \A1[50] , \A1[49] ,
         \A1[48] , \A1[47] , \A1[46] , \A1[45] , \A1[44] , \A1[43] , \A1[42] ,
         \A1[41] , \A1[40] , \A1[39] , \A1[38] , \A1[37] , \A1[36] , \A1[35] ,
         \A1[34] , \A1[33] , \A1[32] , \A1[31] , \A1[30] , \A1[29] , \A1[28] ,
         \A1[27] , \A1[26] , \A1[25] , \A1[24] , \A1[23] , \A1[22] , \A1[21] ,
         \A1[20] , \A1[19] , \A1[18] , \A1[17] , \A1[16] , \A1[15] , \A1[14] ,
         \A1[13] , \A1[12] , \A1[11] , \A1[10] , \A1[9] , \A1[8] , \A1[7] ,
         \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , \A1[1] , \A1[0] ,
         \A2[61] , \A2[60] , \A2[59] , \A2[58] , \A2[57] , \A2[56] , \A2[55] ,
         \A2[54] , \A2[53] , \A2[52] , \A2[51] , \A2[50] , \A2[49] , \A2[48] ,
         \A2[47] , \A2[46] , \A2[45] , \A2[44] , \A2[43] , \A2[42] , \A2[41] ,
         \A2[40] , \A2[39] , \A2[38] , \A2[37] , \A2[36] , \A2[35] , \A2[34] ,
         \A2[33] , \A2[32] , \A2[31] , n4, n5, n6, n7, n8, n9, n10, n11, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28,
         n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42,
         n43, n44, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n57, n58,
         n59, n60, n61, n62, n63, n64, n65, n66, net144709, net144707,
         net144717, net144909, net144973, net145041, net145039, net145037,
         net169226, net169225, net169601, net169776, net169775, net169833,
         \SUMB[31][4] , \SUMB[31][3] , \CARRYB[31][3] , \SUMB[17][15] ,
         \CARRYB[17][15] , \SUMB[30][5] , \SUMB[30][4] , \CARRYB[30][4] ,
         \SUMB[29][6] , \SUMB[29][5] , \CARRYB[29][5] , \SUMB[28][7] ,
         \SUMB[28][6] , \CARRYB[28][6] , \SUMB[27][8] , \SUMB[27][7] ,
         \CARRYB[27][7] , \SUMB[26][9] , \SUMB[26][8] , \CARRYB[26][8] ,
         \SUMB[25][9] , \SUMB[25][10] , \CARRYB[25][9] , \SUMB[24][11] ,
         \SUMB[24][10] , \CARRYB[24][10] , \SUMB[23][12] , \SUMB[23][11] ,
         \CARRYB[23][11] , \SUMB[22][13] , \SUMB[22][12] , \CARRYB[22][12] ,
         \SUMB[21][14] , \SUMB[21][13] , \CARRYB[21][13] , \SUMB[20][15] ,
         \SUMB[20][14] , \CARRYB[20][14] , \SUMB[9][26] , \SUMB[8][27] ,
         \SUMB[7][28] , \SUMB[5][29] , \SUMB[19][16] , \SUMB[19][15] ,
         \SUMB[18][17] , \SUMB[17][18] , \SUMB[16][19] , \SUMB[15][20] ,
         \SUMB[14][21] , \SUMB[13][22] , \SUMB[12][23] , \SUMB[11][24] ,
         \SUMB[10][25] , \CARRYB[9][25] , \CARRYB[8][26] , \CARRYB[7][27] ,
         \CARRYB[6][28] , \CARRYB[19][15] , \CARRYB[18][16] , \CARRYB[17][17] ,
         \CARRYB[16][18] , \CARRYB[15][19] , \CARRYB[14][20] ,
         \CARRYB[13][21] , \CARRYB[12][22] , \CARRYB[11][23] ,
         \CARRYB[10][24] , \SUMB[16][16] , \CARRYB[16][16] , \SUMB[15][17] ,
         \CARRYB[15][17] , \SUMB[14][18] , \CARRYB[14][18] , \SUMB[13][19] ,
         \CARRYB[13][19] , \SUMB[12][20] , \CARRYB[12][20] , \SUMB[11][21] ,
         \CARRYB[11][21] , \SUMB[10][22] , \CARRYB[10][22] , \SUMB[9][23] ,
         \CARRYB[9][23] , \SUMB[8][24] , \CARRYB[8][24] , \SUMB[7][25] ,
         \CARRYB[7][25] , \SUMB[6][26] , \CARRYB[6][26] , \SUMB[5][27] ,
         \CARRYB[5][27] , \SUMB[4][28] , \CARRYB[4][28] , net144713, n56, n45,
         n13, \ab[2][30] , \SUMB[3][29] , \SUMB[2][30] , \CARRYB[3][29] ,
         \CARRYB[2][30] , \SUMB[9][25] , \SUMB[9][24] , \SUMB[8][26] ,
         \SUMB[8][25] , \SUMB[7][27] , \SUMB[7][26] , \SUMB[6][28] ,
         \SUMB[6][27] , \SUMB[5][28] , \SUMB[4][29] , \SUMB[18][16] ,
         \SUMB[18][15] , \SUMB[17][17] , \SUMB[17][16] , \SUMB[16][18] ,
         \SUMB[16][17] , \SUMB[15][19] , \SUMB[15][18] , \SUMB[14][20] ,
         \SUMB[14][19] , \SUMB[13][21] , \SUMB[13][20] , \SUMB[12][22] ,
         \SUMB[12][21] , \SUMB[11][23] , \SUMB[11][22] , \SUMB[10][24] ,
         \SUMB[10][23] , \CARRYB[9][24] , \CARRYB[8][25] , \CARRYB[7][26] ,
         \CARRYB[6][27] , \CARRYB[5][28] , \CARRYB[18][15] , \CARRYB[17][16] ,
         \CARRYB[16][17] , \CARRYB[15][18] , \CARRYB[14][19] ,
         \CARRYB[13][20] , \CARRYB[12][21] , \CARRYB[11][22] ,
         \CARRYB[10][23] , net169827, net169718, net169569, net169256, n67,
         n12, \ab[1][31] , \ab[1][30] , \CARRYB[1][30] , n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102,
         n103, n104, n105, n106, n107, n108, n109, n110, n111, n112, n113,
         n114, n115, n116, n117, n118, n119, n120, n121, n122, n123, n124,
         n125, n126, n127, n128, n129, n130, n131, n132, n133, n134, n135,
         n136, n137, n138, n139, n140, n141, n142, n143, n144, n145, n146,
         n147, n148, n149, n150, n151, n152, n153, n154, n155, n156, n157,
         n158, n159, n160, n161, n162, n163, n164, n165, n166, n167, n168,
         n169, n170, n171, n172, n173, n174, n175, n176, n177, n178, n179,
         n180, n181, n182, n183, n184, n185, n186, n187, n188, n189, n190,
         n191, n192, n193, n194, n195;

  FA_X1 S4_0 ( .A(\ab[31][0] ), .B(\CARRYB[30][0] ), .CI(\SUMB[30][1] ), .CO(
        \CARRYB[31][0] ), .S(\A1[29] ) );
  FA_X1 S4_1 ( .A(\ab[31][1] ), .B(\CARRYB[30][1] ), .CI(\SUMB[30][2] ), .CO(
        \CARRYB[31][1] ), .S(\SUMB[31][1] ) );
  FA_X1 S4_2 ( .A(\ab[31][2] ), .B(\CARRYB[30][2] ), .CI(\SUMB[30][3] ), .CO(
        \CARRYB[31][2] ), .S(\SUMB[31][2] ) );
  FA_X1 S4_5 ( .A(\ab[31][5] ), .B(\CARRYB[30][5] ), .CI(\SUMB[30][6] ), .CO(
        \CARRYB[31][5] ), .S(\SUMB[31][5] ) );
  FA_X1 S4_6 ( .A(\ab[31][6] ), .B(\CARRYB[30][6] ), .CI(\SUMB[30][7] ), .CO(
        \CARRYB[31][6] ), .S(\SUMB[31][6] ) );
  FA_X1 S4_7 ( .A(\ab[31][7] ), .B(\CARRYB[30][7] ), .CI(\SUMB[30][8] ), .CO(
        \CARRYB[31][7] ), .S(\SUMB[31][7] ) );
  FA_X1 S4_8 ( .A(\ab[31][8] ), .B(\CARRYB[30][8] ), .CI(\SUMB[30][9] ), .CO(
        \CARRYB[31][8] ), .S(\SUMB[31][8] ) );
  FA_X1 S4_9 ( .A(\ab[31][9] ), .B(\CARRYB[30][9] ), .CI(\SUMB[30][10] ), .CO(
        \CARRYB[31][9] ), .S(\SUMB[31][9] ) );
  FA_X1 S4_10 ( .A(\ab[31][10] ), .B(\CARRYB[30][10] ), .CI(\SUMB[30][11] ), 
        .CO(\CARRYB[31][10] ), .S(\SUMB[31][10] ) );
  FA_X1 S4_11 ( .A(\ab[31][11] ), .B(\CARRYB[30][11] ), .CI(\SUMB[30][12] ), 
        .CO(\CARRYB[31][11] ), .S(\SUMB[31][11] ) );
  FA_X1 S4_12 ( .A(\ab[31][12] ), .B(\CARRYB[30][12] ), .CI(\SUMB[30][13] ), 
        .CO(\CARRYB[31][12] ), .S(\SUMB[31][12] ) );
  FA_X1 S4_13 ( .A(\ab[31][13] ), .B(\CARRYB[30][13] ), .CI(\SUMB[30][14] ), 
        .CO(\CARRYB[31][13] ), .S(\SUMB[31][13] ) );
  FA_X1 S4_14 ( .A(\ab[31][14] ), .B(\CARRYB[30][14] ), .CI(\SUMB[30][15] ), 
        .CO(\CARRYB[31][14] ), .S(\SUMB[31][14] ) );
  FA_X1 S4_15 ( .A(\ab[31][15] ), .B(\CARRYB[30][15] ), .CI(\SUMB[30][16] ), 
        .CO(\CARRYB[31][15] ), .S(\SUMB[31][15] ) );
  FA_X1 S4_16 ( .A(\ab[31][16] ), .B(\CARRYB[30][16] ), .CI(\SUMB[30][17] ), 
        .CO(\CARRYB[31][16] ), .S(\SUMB[31][16] ) );
  FA_X1 S4_17 ( .A(\ab[31][17] ), .B(\CARRYB[30][17] ), .CI(\SUMB[30][18] ), 
        .CO(\CARRYB[31][17] ), .S(\SUMB[31][17] ) );
  FA_X1 S4_18 ( .A(\ab[31][18] ), .B(\CARRYB[30][18] ), .CI(\SUMB[30][19] ), 
        .CO(\CARRYB[31][18] ), .S(\SUMB[31][18] ) );
  FA_X1 S4_19 ( .A(\ab[31][19] ), .B(\CARRYB[30][19] ), .CI(\SUMB[30][20] ), 
        .CO(\CARRYB[31][19] ), .S(\SUMB[31][19] ) );
  FA_X1 S4_20 ( .A(\ab[31][20] ), .B(\CARRYB[30][20] ), .CI(\SUMB[30][21] ), 
        .CO(\CARRYB[31][20] ), .S(\SUMB[31][20] ) );
  FA_X1 S4_21 ( .A(\ab[31][21] ), .B(\CARRYB[30][21] ), .CI(\SUMB[30][22] ), 
        .CO(\CARRYB[31][21] ), .S(\SUMB[31][21] ) );
  FA_X1 S4_22 ( .A(\ab[31][22] ), .B(\CARRYB[30][22] ), .CI(\SUMB[30][23] ), 
        .CO(\CARRYB[31][22] ), .S(\SUMB[31][22] ) );
  FA_X1 S4_23 ( .A(\ab[31][23] ), .B(\CARRYB[30][23] ), .CI(\SUMB[30][24] ), 
        .CO(\CARRYB[31][23] ), .S(\SUMB[31][23] ) );
  FA_X1 S4_24 ( .A(\ab[31][24] ), .B(\CARRYB[30][24] ), .CI(\SUMB[30][25] ), 
        .CO(\CARRYB[31][24] ), .S(\SUMB[31][24] ) );
  FA_X1 S4_25 ( .A(\ab[31][25] ), .B(\CARRYB[30][25] ), .CI(\SUMB[30][26] ), 
        .CO(\CARRYB[31][25] ), .S(\SUMB[31][25] ) );
  FA_X1 S4_26 ( .A(\ab[31][26] ), .B(\CARRYB[30][26] ), .CI(\SUMB[30][27] ), 
        .CO(\CARRYB[31][26] ), .S(\SUMB[31][26] ) );
  FA_X1 S4_27 ( .A(\ab[31][27] ), .B(\CARRYB[30][27] ), .CI(\SUMB[30][28] ), 
        .CO(\CARRYB[31][27] ), .S(\SUMB[31][27] ) );
  FA_X1 S4_28 ( .A(\ab[31][28] ), .B(\CARRYB[30][28] ), .CI(\SUMB[30][29] ), 
        .CO(\CARRYB[31][28] ), .S(\SUMB[31][28] ) );
  FA_X1 S4_29 ( .A(\ab[31][29] ), .B(\CARRYB[30][29] ), .CI(\SUMB[30][30] ), 
        .CO(\CARRYB[31][29] ), .S(\SUMB[31][29] ) );
  FA_X1 S5_30 ( .A(\ab[31][30] ), .B(\CARRYB[30][30] ), .CI(\ab[30][31] ), 
        .CO(\CARRYB[31][30] ), .S(\SUMB[31][30] ) );
  FA_X1 S1_30_0 ( .A(\ab[30][0] ), .B(\CARRYB[29][0] ), .CI(\SUMB[29][1] ), 
        .CO(\CARRYB[30][0] ), .S(\A1[28] ) );
  FA_X1 S2_30_1 ( .A(\ab[30][1] ), .B(\CARRYB[29][1] ), .CI(\SUMB[29][2] ), 
        .CO(\CARRYB[30][1] ), .S(\SUMB[30][1] ) );
  FA_X1 S2_30_2 ( .A(\ab[30][2] ), .B(\CARRYB[29][2] ), .CI(\SUMB[29][3] ), 
        .CO(\CARRYB[30][2] ), .S(\SUMB[30][2] ) );
  FA_X1 S2_30_3 ( .A(\CARRYB[29][3] ), .B(\ab[30][3] ), .CI(\SUMB[29][4] ), 
        .CO(\CARRYB[30][3] ), .S(\SUMB[30][3] ) );
  FA_X1 S2_30_6 ( .A(\ab[30][6] ), .B(\CARRYB[29][6] ), .CI(\SUMB[29][7] ), 
        .CO(\CARRYB[30][6] ), .S(\SUMB[30][6] ) );
  FA_X1 S2_30_7 ( .A(\ab[30][7] ), .B(\CARRYB[29][7] ), .CI(\SUMB[29][8] ), 
        .CO(\CARRYB[30][7] ), .S(\SUMB[30][7] ) );
  FA_X1 S2_30_8 ( .A(\ab[30][8] ), .B(\CARRYB[29][8] ), .CI(\SUMB[29][9] ), 
        .CO(\CARRYB[30][8] ), .S(\SUMB[30][8] ) );
  FA_X1 S2_30_9 ( .A(\ab[30][9] ), .B(\CARRYB[29][9] ), .CI(\SUMB[29][10] ), 
        .CO(\CARRYB[30][9] ), .S(\SUMB[30][9] ) );
  FA_X1 S2_30_10 ( .A(\ab[30][10] ), .B(\CARRYB[29][10] ), .CI(\SUMB[29][11] ), 
        .CO(\CARRYB[30][10] ), .S(\SUMB[30][10] ) );
  FA_X1 S2_30_11 ( .A(\ab[30][11] ), .B(\CARRYB[29][11] ), .CI(\SUMB[29][12] ), 
        .CO(\CARRYB[30][11] ), .S(\SUMB[30][11] ) );
  FA_X1 S2_30_12 ( .A(\ab[30][12] ), .B(\CARRYB[29][12] ), .CI(\SUMB[29][13] ), 
        .CO(\CARRYB[30][12] ), .S(\SUMB[30][12] ) );
  FA_X1 S2_30_13 ( .A(\ab[30][13] ), .B(\CARRYB[29][13] ), .CI(\SUMB[29][14] ), 
        .CO(\CARRYB[30][13] ), .S(\SUMB[30][13] ) );
  FA_X1 S2_30_14 ( .A(\ab[30][14] ), .B(\CARRYB[29][14] ), .CI(\SUMB[29][15] ), 
        .CO(\CARRYB[30][14] ), .S(\SUMB[30][14] ) );
  FA_X1 S2_30_15 ( .A(\ab[30][15] ), .B(\CARRYB[29][15] ), .CI(\SUMB[29][16] ), 
        .CO(\CARRYB[30][15] ), .S(\SUMB[30][15] ) );
  FA_X1 S2_30_16 ( .A(\ab[30][16] ), .B(\CARRYB[29][16] ), .CI(\SUMB[29][17] ), 
        .CO(\CARRYB[30][16] ), .S(\SUMB[30][16] ) );
  FA_X1 S2_30_17 ( .A(\ab[30][17] ), .B(\CARRYB[29][17] ), .CI(\SUMB[29][18] ), 
        .CO(\CARRYB[30][17] ), .S(\SUMB[30][17] ) );
  FA_X1 S2_30_18 ( .A(\ab[30][18] ), .B(\CARRYB[29][18] ), .CI(\SUMB[29][19] ), 
        .CO(\CARRYB[30][18] ), .S(\SUMB[30][18] ) );
  FA_X1 S2_30_19 ( .A(\ab[30][19] ), .B(\CARRYB[29][19] ), .CI(\SUMB[29][20] ), 
        .CO(\CARRYB[30][19] ), .S(\SUMB[30][19] ) );
  FA_X1 S2_30_20 ( .A(\ab[30][20] ), .B(\CARRYB[29][20] ), .CI(\SUMB[29][21] ), 
        .CO(\CARRYB[30][20] ), .S(\SUMB[30][20] ) );
  FA_X1 S2_30_21 ( .A(\ab[30][21] ), .B(\CARRYB[29][21] ), .CI(\SUMB[29][22] ), 
        .CO(\CARRYB[30][21] ), .S(\SUMB[30][21] ) );
  FA_X1 S2_30_22 ( .A(\ab[30][22] ), .B(\CARRYB[29][22] ), .CI(\SUMB[29][23] ), 
        .CO(\CARRYB[30][22] ), .S(\SUMB[30][22] ) );
  FA_X1 S2_30_23 ( .A(\ab[30][23] ), .B(\CARRYB[29][23] ), .CI(\SUMB[29][24] ), 
        .CO(\CARRYB[30][23] ), .S(\SUMB[30][23] ) );
  FA_X1 S2_30_24 ( .A(\ab[30][24] ), .B(\CARRYB[29][24] ), .CI(\SUMB[29][25] ), 
        .CO(\CARRYB[30][24] ), .S(\SUMB[30][24] ) );
  FA_X1 S2_30_25 ( .A(\ab[30][25] ), .B(\CARRYB[29][25] ), .CI(\SUMB[29][26] ), 
        .CO(\CARRYB[30][25] ), .S(\SUMB[30][25] ) );
  FA_X1 S2_30_26 ( .A(\ab[30][26] ), .B(\CARRYB[29][26] ), .CI(\SUMB[29][27] ), 
        .CO(\CARRYB[30][26] ), .S(\SUMB[30][26] ) );
  FA_X1 S2_30_27 ( .A(\ab[30][27] ), .B(\CARRYB[29][27] ), .CI(\SUMB[29][28] ), 
        .CO(\CARRYB[30][27] ), .S(\SUMB[30][27] ) );
  FA_X1 S2_30_28 ( .A(\ab[30][28] ), .B(\CARRYB[29][28] ), .CI(\SUMB[29][29] ), 
        .CO(\CARRYB[30][28] ), .S(\SUMB[30][28] ) );
  FA_X1 S2_30_29 ( .A(\ab[30][29] ), .B(\CARRYB[29][29] ), .CI(\SUMB[29][30] ), 
        .CO(\CARRYB[30][29] ), .S(\SUMB[30][29] ) );
  FA_X1 S3_30_30 ( .A(\ab[30][30] ), .B(\CARRYB[29][30] ), .CI(\ab[29][31] ), 
        .CO(\CARRYB[30][30] ), .S(\SUMB[30][30] ) );
  FA_X1 S1_29_0 ( .A(\ab[29][0] ), .B(\CARRYB[28][0] ), .CI(\SUMB[28][1] ), 
        .CO(\CARRYB[29][0] ), .S(\A1[27] ) );
  FA_X1 S2_29_1 ( .A(\ab[29][1] ), .B(\CARRYB[28][1] ), .CI(\SUMB[28][2] ), 
        .CO(\CARRYB[29][1] ), .S(\SUMB[29][1] ) );
  FA_X1 S2_29_2 ( .A(\ab[29][2] ), .B(\CARRYB[28][2] ), .CI(\SUMB[28][3] ), 
        .CO(\CARRYB[29][2] ), .S(\SUMB[29][2] ) );
  FA_X1 S2_29_3 ( .A(\CARRYB[28][3] ), .B(\ab[29][3] ), .CI(\SUMB[28][4] ), 
        .CO(\CARRYB[29][3] ), .S(\SUMB[29][3] ) );
  FA_X1 S2_29_4 ( .A(\ab[29][4] ), .B(\CARRYB[28][4] ), .CI(\SUMB[28][5] ), 
        .CO(\CARRYB[29][4] ), .S(\SUMB[29][4] ) );
  FA_X1 S2_29_7 ( .A(\ab[29][7] ), .B(\CARRYB[28][7] ), .CI(\SUMB[28][8] ), 
        .CO(\CARRYB[29][7] ), .S(\SUMB[29][7] ) );
  FA_X1 S2_29_8 ( .A(\ab[29][8] ), .B(\CARRYB[28][8] ), .CI(\SUMB[28][9] ), 
        .CO(\CARRYB[29][8] ), .S(\SUMB[29][8] ) );
  FA_X1 S2_29_9 ( .A(\ab[29][9] ), .B(\CARRYB[28][9] ), .CI(\SUMB[28][10] ), 
        .CO(\CARRYB[29][9] ), .S(\SUMB[29][9] ) );
  FA_X1 S2_29_10 ( .A(\ab[29][10] ), .B(\CARRYB[28][10] ), .CI(\SUMB[28][11] ), 
        .CO(\CARRYB[29][10] ), .S(\SUMB[29][10] ) );
  FA_X1 S2_29_11 ( .A(\ab[29][11] ), .B(\CARRYB[28][11] ), .CI(\SUMB[28][12] ), 
        .CO(\CARRYB[29][11] ), .S(\SUMB[29][11] ) );
  FA_X1 S2_29_12 ( .A(\ab[29][12] ), .B(\CARRYB[28][12] ), .CI(\SUMB[28][13] ), 
        .CO(\CARRYB[29][12] ), .S(\SUMB[29][12] ) );
  FA_X1 S2_29_13 ( .A(\ab[29][13] ), .B(\CARRYB[28][13] ), .CI(\SUMB[28][14] ), 
        .CO(\CARRYB[29][13] ), .S(\SUMB[29][13] ) );
  FA_X1 S2_29_14 ( .A(\ab[29][14] ), .B(\CARRYB[28][14] ), .CI(\SUMB[28][15] ), 
        .CO(\CARRYB[29][14] ), .S(\SUMB[29][14] ) );
  FA_X1 S2_29_15 ( .A(\ab[29][15] ), .B(\CARRYB[28][15] ), .CI(\SUMB[28][16] ), 
        .CO(\CARRYB[29][15] ), .S(\SUMB[29][15] ) );
  FA_X1 S2_29_16 ( .A(\ab[29][16] ), .B(\CARRYB[28][16] ), .CI(\SUMB[28][17] ), 
        .CO(\CARRYB[29][16] ), .S(\SUMB[29][16] ) );
  FA_X1 S2_29_17 ( .A(\ab[29][17] ), .B(\CARRYB[28][17] ), .CI(\SUMB[28][18] ), 
        .CO(\CARRYB[29][17] ), .S(\SUMB[29][17] ) );
  FA_X1 S2_29_18 ( .A(\ab[29][18] ), .B(\CARRYB[28][18] ), .CI(\SUMB[28][19] ), 
        .CO(\CARRYB[29][18] ), .S(\SUMB[29][18] ) );
  FA_X1 S2_29_19 ( .A(\ab[29][19] ), .B(\CARRYB[28][19] ), .CI(\SUMB[28][20] ), 
        .CO(\CARRYB[29][19] ), .S(\SUMB[29][19] ) );
  FA_X1 S2_29_20 ( .A(\ab[29][20] ), .B(\CARRYB[28][20] ), .CI(\SUMB[28][21] ), 
        .CO(\CARRYB[29][20] ), .S(\SUMB[29][20] ) );
  FA_X1 S2_29_21 ( .A(\ab[29][21] ), .B(\CARRYB[28][21] ), .CI(\SUMB[28][22] ), 
        .CO(\CARRYB[29][21] ), .S(\SUMB[29][21] ) );
  FA_X1 S2_29_22 ( .A(\ab[29][22] ), .B(\CARRYB[28][22] ), .CI(\SUMB[28][23] ), 
        .CO(\CARRYB[29][22] ), .S(\SUMB[29][22] ) );
  FA_X1 S2_29_23 ( .A(\ab[29][23] ), .B(\CARRYB[28][23] ), .CI(\SUMB[28][24] ), 
        .CO(\CARRYB[29][23] ), .S(\SUMB[29][23] ) );
  FA_X1 S2_29_24 ( .A(\ab[29][24] ), .B(\CARRYB[28][24] ), .CI(\SUMB[28][25] ), 
        .CO(\CARRYB[29][24] ), .S(\SUMB[29][24] ) );
  FA_X1 S2_29_25 ( .A(\ab[29][25] ), .B(\CARRYB[28][25] ), .CI(\SUMB[28][26] ), 
        .CO(\CARRYB[29][25] ), .S(\SUMB[29][25] ) );
  FA_X1 S2_29_26 ( .A(\ab[29][26] ), .B(\CARRYB[28][26] ), .CI(\SUMB[28][27] ), 
        .CO(\CARRYB[29][26] ), .S(\SUMB[29][26] ) );
  FA_X1 S2_29_27 ( .A(\ab[29][27] ), .B(\CARRYB[28][27] ), .CI(\SUMB[28][28] ), 
        .CO(\CARRYB[29][27] ), .S(\SUMB[29][27] ) );
  FA_X1 S2_29_28 ( .A(\ab[29][28] ), .B(\CARRYB[28][28] ), .CI(\SUMB[28][29] ), 
        .CO(\CARRYB[29][28] ), .S(\SUMB[29][28] ) );
  FA_X1 S2_29_29 ( .A(\ab[29][29] ), .B(\CARRYB[28][29] ), .CI(\SUMB[28][30] ), 
        .CO(\CARRYB[29][29] ), .S(\SUMB[29][29] ) );
  FA_X1 S3_29_30 ( .A(\ab[29][30] ), .B(\CARRYB[28][30] ), .CI(\ab[28][31] ), 
        .CO(\CARRYB[29][30] ), .S(\SUMB[29][30] ) );
  FA_X1 S1_28_0 ( .A(\ab[28][0] ), .B(\CARRYB[27][0] ), .CI(\SUMB[27][1] ), 
        .CO(\CARRYB[28][0] ), .S(\A1[26] ) );
  FA_X1 S2_28_1 ( .A(\ab[28][1] ), .B(\CARRYB[27][1] ), .CI(\SUMB[27][2] ), 
        .CO(\CARRYB[28][1] ), .S(\SUMB[28][1] ) );
  FA_X1 S2_28_2 ( .A(\ab[28][2] ), .B(\CARRYB[27][2] ), .CI(\SUMB[27][3] ), 
        .CO(\CARRYB[28][2] ), .S(\SUMB[28][2] ) );
  FA_X1 S2_28_3 ( .A(\ab[28][3] ), .B(\CARRYB[27][3] ), .CI(\SUMB[27][4] ), 
        .CO(\CARRYB[28][3] ), .S(\SUMB[28][3] ) );
  FA_X1 S2_28_4 ( .A(\ab[28][4] ), .B(\CARRYB[27][4] ), .CI(\SUMB[27][5] ), 
        .CO(\CARRYB[28][4] ), .S(\SUMB[28][4] ) );
  FA_X1 S2_28_5 ( .A(\CARRYB[27][5] ), .B(\ab[28][5] ), .CI(\SUMB[27][6] ), 
        .CO(\CARRYB[28][5] ), .S(\SUMB[28][5] ) );
  FA_X1 S2_28_8 ( .A(\ab[28][8] ), .B(\CARRYB[27][8] ), .CI(\SUMB[27][9] ), 
        .CO(\CARRYB[28][8] ), .S(\SUMB[28][8] ) );
  FA_X1 S2_28_9 ( .A(\ab[28][9] ), .B(\CARRYB[27][9] ), .CI(\SUMB[27][10] ), 
        .CO(\CARRYB[28][9] ), .S(\SUMB[28][9] ) );
  FA_X1 S2_28_10 ( .A(\ab[28][10] ), .B(\CARRYB[27][10] ), .CI(\SUMB[27][11] ), 
        .CO(\CARRYB[28][10] ), .S(\SUMB[28][10] ) );
  FA_X1 S2_28_11 ( .A(\ab[28][11] ), .B(\CARRYB[27][11] ), .CI(\SUMB[27][12] ), 
        .CO(\CARRYB[28][11] ), .S(\SUMB[28][11] ) );
  FA_X1 S2_28_12 ( .A(\ab[28][12] ), .B(\CARRYB[27][12] ), .CI(\SUMB[27][13] ), 
        .CO(\CARRYB[28][12] ), .S(\SUMB[28][12] ) );
  FA_X1 S2_28_13 ( .A(\ab[28][13] ), .B(\CARRYB[27][13] ), .CI(\SUMB[27][14] ), 
        .CO(\CARRYB[28][13] ), .S(\SUMB[28][13] ) );
  FA_X1 S2_28_14 ( .A(\ab[28][14] ), .B(\CARRYB[27][14] ), .CI(\SUMB[27][15] ), 
        .CO(\CARRYB[28][14] ), .S(\SUMB[28][14] ) );
  FA_X1 S2_28_15 ( .A(\ab[28][15] ), .B(\CARRYB[27][15] ), .CI(\SUMB[27][16] ), 
        .CO(\CARRYB[28][15] ), .S(\SUMB[28][15] ) );
  FA_X1 S2_28_16 ( .A(\ab[28][16] ), .B(\CARRYB[27][16] ), .CI(\SUMB[27][17] ), 
        .CO(\CARRYB[28][16] ), .S(\SUMB[28][16] ) );
  FA_X1 S2_28_17 ( .A(\ab[28][17] ), .B(\CARRYB[27][17] ), .CI(\SUMB[27][18] ), 
        .CO(\CARRYB[28][17] ), .S(\SUMB[28][17] ) );
  FA_X1 S2_28_18 ( .A(\ab[28][18] ), .B(\CARRYB[27][18] ), .CI(\SUMB[27][19] ), 
        .CO(\CARRYB[28][18] ), .S(\SUMB[28][18] ) );
  FA_X1 S2_28_19 ( .A(\ab[28][19] ), .B(\CARRYB[27][19] ), .CI(\SUMB[27][20] ), 
        .CO(\CARRYB[28][19] ), .S(\SUMB[28][19] ) );
  FA_X1 S2_28_20 ( .A(\ab[28][20] ), .B(\CARRYB[27][20] ), .CI(\SUMB[27][21] ), 
        .CO(\CARRYB[28][20] ), .S(\SUMB[28][20] ) );
  FA_X1 S2_28_21 ( .A(\ab[28][21] ), .B(\CARRYB[27][21] ), .CI(\SUMB[27][22] ), 
        .CO(\CARRYB[28][21] ), .S(\SUMB[28][21] ) );
  FA_X1 S2_28_22 ( .A(\ab[28][22] ), .B(\CARRYB[27][22] ), .CI(\SUMB[27][23] ), 
        .CO(\CARRYB[28][22] ), .S(\SUMB[28][22] ) );
  FA_X1 S2_28_23 ( .A(\ab[28][23] ), .B(\CARRYB[27][23] ), .CI(\SUMB[27][24] ), 
        .CO(\CARRYB[28][23] ), .S(\SUMB[28][23] ) );
  FA_X1 S2_28_24 ( .A(\ab[28][24] ), .B(\CARRYB[27][24] ), .CI(\SUMB[27][25] ), 
        .CO(\CARRYB[28][24] ), .S(\SUMB[28][24] ) );
  FA_X1 S2_28_25 ( .A(\ab[28][25] ), .B(\CARRYB[27][25] ), .CI(\SUMB[27][26] ), 
        .CO(\CARRYB[28][25] ), .S(\SUMB[28][25] ) );
  FA_X1 S2_28_26 ( .A(\ab[28][26] ), .B(\CARRYB[27][26] ), .CI(\SUMB[27][27] ), 
        .CO(\CARRYB[28][26] ), .S(\SUMB[28][26] ) );
  FA_X1 S2_28_27 ( .A(\ab[28][27] ), .B(\CARRYB[27][27] ), .CI(\SUMB[27][28] ), 
        .CO(\CARRYB[28][27] ), .S(\SUMB[28][27] ) );
  FA_X1 S2_28_28 ( .A(\ab[28][28] ), .B(\CARRYB[27][28] ), .CI(\SUMB[27][29] ), 
        .CO(\CARRYB[28][28] ), .S(\SUMB[28][28] ) );
  FA_X1 S2_28_29 ( .A(\ab[28][29] ), .B(\CARRYB[27][29] ), .CI(\SUMB[27][30] ), 
        .CO(\CARRYB[28][29] ), .S(\SUMB[28][29] ) );
  FA_X1 S3_28_30 ( .A(\ab[28][30] ), .B(\CARRYB[27][30] ), .CI(\ab[27][31] ), 
        .CO(\CARRYB[28][30] ), .S(\SUMB[28][30] ) );
  FA_X1 S1_27_0 ( .A(\ab[27][0] ), .B(\CARRYB[26][0] ), .CI(\SUMB[26][1] ), 
        .CO(\CARRYB[27][0] ), .S(\A1[25] ) );
  FA_X1 S2_27_1 ( .A(\ab[27][1] ), .B(\CARRYB[26][1] ), .CI(\SUMB[26][2] ), 
        .CO(\CARRYB[27][1] ), .S(\SUMB[27][1] ) );
  FA_X1 S2_27_2 ( .A(\ab[27][2] ), .B(\CARRYB[26][2] ), .CI(\SUMB[26][3] ), 
        .CO(\CARRYB[27][2] ), .S(\SUMB[27][2] ) );
  FA_X1 S2_27_3 ( .A(\ab[27][3] ), .B(\CARRYB[26][3] ), .CI(\SUMB[26][4] ), 
        .CO(\CARRYB[27][3] ), .S(\SUMB[27][3] ) );
  FA_X1 S2_27_4 ( .A(\ab[27][4] ), .B(\CARRYB[26][4] ), .CI(\SUMB[26][5] ), 
        .CO(\CARRYB[27][4] ), .S(\SUMB[27][4] ) );
  FA_X1 S2_27_5 ( .A(\CARRYB[26][5] ), .B(\ab[27][5] ), .CI(\SUMB[26][6] ), 
        .CO(\CARRYB[27][5] ), .S(\SUMB[27][5] ) );
  FA_X1 S2_27_6 ( .A(\ab[27][6] ), .B(\CARRYB[26][6] ), .CI(\SUMB[26][7] ), 
        .CO(\CARRYB[27][6] ), .S(\SUMB[27][6] ) );
  FA_X1 S2_27_9 ( .A(\ab[27][9] ), .B(\CARRYB[26][9] ), .CI(\SUMB[26][10] ), 
        .CO(\CARRYB[27][9] ), .S(\SUMB[27][9] ) );
  FA_X1 S2_27_10 ( .A(\ab[27][10] ), .B(\CARRYB[26][10] ), .CI(\SUMB[26][11] ), 
        .CO(\CARRYB[27][10] ), .S(\SUMB[27][10] ) );
  FA_X1 S2_27_11 ( .A(\ab[27][11] ), .B(\CARRYB[26][11] ), .CI(\SUMB[26][12] ), 
        .CO(\CARRYB[27][11] ), .S(\SUMB[27][11] ) );
  FA_X1 S2_27_12 ( .A(\ab[27][12] ), .B(\CARRYB[26][12] ), .CI(\SUMB[26][13] ), 
        .CO(\CARRYB[27][12] ), .S(\SUMB[27][12] ) );
  FA_X1 S2_27_13 ( .A(\ab[27][13] ), .B(\CARRYB[26][13] ), .CI(\SUMB[26][14] ), 
        .CO(\CARRYB[27][13] ), .S(\SUMB[27][13] ) );
  FA_X1 S2_27_14 ( .A(\ab[27][14] ), .B(\CARRYB[26][14] ), .CI(\SUMB[26][15] ), 
        .CO(\CARRYB[27][14] ), .S(\SUMB[27][14] ) );
  FA_X1 S2_27_15 ( .A(\ab[27][15] ), .B(\CARRYB[26][15] ), .CI(\SUMB[26][16] ), 
        .CO(\CARRYB[27][15] ), .S(\SUMB[27][15] ) );
  FA_X1 S2_27_16 ( .A(\ab[27][16] ), .B(\CARRYB[26][16] ), .CI(\SUMB[26][17] ), 
        .CO(\CARRYB[27][16] ), .S(\SUMB[27][16] ) );
  FA_X1 S2_27_17 ( .A(\ab[27][17] ), .B(\CARRYB[26][17] ), .CI(\SUMB[26][18] ), 
        .CO(\CARRYB[27][17] ), .S(\SUMB[27][17] ) );
  FA_X1 S2_27_18 ( .A(\ab[27][18] ), .B(\CARRYB[26][18] ), .CI(\SUMB[26][19] ), 
        .CO(\CARRYB[27][18] ), .S(\SUMB[27][18] ) );
  FA_X1 S2_27_19 ( .A(\ab[27][19] ), .B(\CARRYB[26][19] ), .CI(\SUMB[26][20] ), 
        .CO(\CARRYB[27][19] ), .S(\SUMB[27][19] ) );
  FA_X1 S2_27_20 ( .A(\ab[27][20] ), .B(\CARRYB[26][20] ), .CI(\SUMB[26][21] ), 
        .CO(\CARRYB[27][20] ), .S(\SUMB[27][20] ) );
  FA_X1 S2_27_21 ( .A(\ab[27][21] ), .B(\CARRYB[26][21] ), .CI(\SUMB[26][22] ), 
        .CO(\CARRYB[27][21] ), .S(\SUMB[27][21] ) );
  FA_X1 S2_27_22 ( .A(\ab[27][22] ), .B(\CARRYB[26][22] ), .CI(\SUMB[26][23] ), 
        .CO(\CARRYB[27][22] ), .S(\SUMB[27][22] ) );
  FA_X1 S2_27_23 ( .A(\ab[27][23] ), .B(\CARRYB[26][23] ), .CI(\SUMB[26][24] ), 
        .CO(\CARRYB[27][23] ), .S(\SUMB[27][23] ) );
  FA_X1 S2_27_24 ( .A(\ab[27][24] ), .B(\CARRYB[26][24] ), .CI(\SUMB[26][25] ), 
        .CO(\CARRYB[27][24] ), .S(\SUMB[27][24] ) );
  FA_X1 S2_27_25 ( .A(\ab[27][25] ), .B(\CARRYB[26][25] ), .CI(\SUMB[26][26] ), 
        .CO(\CARRYB[27][25] ), .S(\SUMB[27][25] ) );
  FA_X1 S2_27_26 ( .A(\ab[27][26] ), .B(\CARRYB[26][26] ), .CI(\SUMB[26][27] ), 
        .CO(\CARRYB[27][26] ), .S(\SUMB[27][26] ) );
  FA_X1 S2_27_27 ( .A(\ab[27][27] ), .B(\CARRYB[26][27] ), .CI(\SUMB[26][28] ), 
        .CO(\CARRYB[27][27] ), .S(\SUMB[27][27] ) );
  FA_X1 S2_27_28 ( .A(\ab[27][28] ), .B(\CARRYB[26][28] ), .CI(\SUMB[26][29] ), 
        .CO(\CARRYB[27][28] ), .S(\SUMB[27][28] ) );
  FA_X1 S2_27_29 ( .A(\ab[27][29] ), .B(\CARRYB[26][29] ), .CI(\SUMB[26][30] ), 
        .CO(\CARRYB[27][29] ), .S(\SUMB[27][29] ) );
  FA_X1 S3_27_30 ( .A(\ab[27][30] ), .B(\CARRYB[26][30] ), .CI(\ab[26][31] ), 
        .CO(\CARRYB[27][30] ), .S(\SUMB[27][30] ) );
  FA_X1 S1_26_0 ( .A(\ab[26][0] ), .B(\CARRYB[25][0] ), .CI(\SUMB[25][1] ), 
        .CO(\CARRYB[26][0] ), .S(\A1[24] ) );
  FA_X1 S2_26_1 ( .A(\ab[26][1] ), .B(\CARRYB[25][1] ), .CI(\SUMB[25][2] ), 
        .CO(\CARRYB[26][1] ), .S(\SUMB[26][1] ) );
  FA_X1 S2_26_2 ( .A(\ab[26][2] ), .B(\CARRYB[25][2] ), .CI(\SUMB[25][3] ), 
        .CO(\CARRYB[26][2] ), .S(\SUMB[26][2] ) );
  FA_X1 S2_26_3 ( .A(\ab[26][3] ), .B(\CARRYB[25][3] ), .CI(\SUMB[25][4] ), 
        .CO(\CARRYB[26][3] ), .S(\SUMB[26][3] ) );
  FA_X1 S2_26_4 ( .A(\ab[26][4] ), .B(\CARRYB[25][4] ), .CI(\SUMB[25][5] ), 
        .CO(\CARRYB[26][4] ), .S(\SUMB[26][4] ) );
  FA_X1 S2_26_5 ( .A(\ab[26][5] ), .B(\CARRYB[25][5] ), .CI(\SUMB[25][6] ), 
        .CO(\CARRYB[26][5] ), .S(\SUMB[26][5] ) );
  FA_X1 S2_26_6 ( .A(\ab[26][6] ), .B(\CARRYB[25][6] ), .CI(\SUMB[25][7] ), 
        .CO(\CARRYB[26][6] ), .S(\SUMB[26][6] ) );
  FA_X1 S2_26_7 ( .A(\CARRYB[25][7] ), .B(\ab[26][7] ), .CI(\SUMB[25][8] ), 
        .CO(\CARRYB[26][7] ), .S(\SUMB[26][7] ) );
  FA_X1 S2_26_10 ( .A(\ab[26][10] ), .B(\CARRYB[25][10] ), .CI(\SUMB[25][11] ), 
        .CO(\CARRYB[26][10] ), .S(\SUMB[26][10] ) );
  FA_X1 S2_26_11 ( .A(\ab[26][11] ), .B(\CARRYB[25][11] ), .CI(\SUMB[25][12] ), 
        .CO(\CARRYB[26][11] ), .S(\SUMB[26][11] ) );
  FA_X1 S2_26_12 ( .A(\ab[26][12] ), .B(\CARRYB[25][12] ), .CI(\SUMB[25][13] ), 
        .CO(\CARRYB[26][12] ), .S(\SUMB[26][12] ) );
  FA_X1 S2_26_13 ( .A(\ab[26][13] ), .B(\CARRYB[25][13] ), .CI(\SUMB[25][14] ), 
        .CO(\CARRYB[26][13] ), .S(\SUMB[26][13] ) );
  FA_X1 S2_26_14 ( .A(\ab[26][14] ), .B(\CARRYB[25][14] ), .CI(\SUMB[25][15] ), 
        .CO(\CARRYB[26][14] ), .S(\SUMB[26][14] ) );
  FA_X1 S2_26_15 ( .A(\ab[26][15] ), .B(\CARRYB[25][15] ), .CI(\SUMB[25][16] ), 
        .CO(\CARRYB[26][15] ), .S(\SUMB[26][15] ) );
  FA_X1 S2_26_16 ( .A(\ab[26][16] ), .B(\CARRYB[25][16] ), .CI(\SUMB[25][17] ), 
        .CO(\CARRYB[26][16] ), .S(\SUMB[26][16] ) );
  FA_X1 S2_26_17 ( .A(\ab[26][17] ), .B(\CARRYB[25][17] ), .CI(\SUMB[25][18] ), 
        .CO(\CARRYB[26][17] ), .S(\SUMB[26][17] ) );
  FA_X1 S2_26_18 ( .A(\ab[26][18] ), .B(\CARRYB[25][18] ), .CI(\SUMB[25][19] ), 
        .CO(\CARRYB[26][18] ), .S(\SUMB[26][18] ) );
  FA_X1 S2_26_19 ( .A(\ab[26][19] ), .B(\CARRYB[25][19] ), .CI(\SUMB[25][20] ), 
        .CO(\CARRYB[26][19] ), .S(\SUMB[26][19] ) );
  FA_X1 S2_26_20 ( .A(\ab[26][20] ), .B(\CARRYB[25][20] ), .CI(\SUMB[25][21] ), 
        .CO(\CARRYB[26][20] ), .S(\SUMB[26][20] ) );
  FA_X1 S2_26_21 ( .A(\ab[26][21] ), .B(\CARRYB[25][21] ), .CI(\SUMB[25][22] ), 
        .CO(\CARRYB[26][21] ), .S(\SUMB[26][21] ) );
  FA_X1 S2_26_22 ( .A(\ab[26][22] ), .B(\CARRYB[25][22] ), .CI(\SUMB[25][23] ), 
        .CO(\CARRYB[26][22] ), .S(\SUMB[26][22] ) );
  FA_X1 S2_26_23 ( .A(\ab[26][23] ), .B(\CARRYB[25][23] ), .CI(\SUMB[25][24] ), 
        .CO(\CARRYB[26][23] ), .S(\SUMB[26][23] ) );
  FA_X1 S2_26_24 ( .A(\ab[26][24] ), .B(\CARRYB[25][24] ), .CI(\SUMB[25][25] ), 
        .CO(\CARRYB[26][24] ), .S(\SUMB[26][24] ) );
  FA_X1 S2_26_25 ( .A(\ab[26][25] ), .B(\CARRYB[25][25] ), .CI(\SUMB[25][26] ), 
        .CO(\CARRYB[26][25] ), .S(\SUMB[26][25] ) );
  FA_X1 S2_26_26 ( .A(\ab[26][26] ), .B(\CARRYB[25][26] ), .CI(\SUMB[25][27] ), 
        .CO(\CARRYB[26][26] ), .S(\SUMB[26][26] ) );
  FA_X1 S2_26_27 ( .A(\ab[26][27] ), .B(\CARRYB[25][27] ), .CI(\SUMB[25][28] ), 
        .CO(\CARRYB[26][27] ), .S(\SUMB[26][27] ) );
  FA_X1 S2_26_28 ( .A(\ab[26][28] ), .B(\CARRYB[25][28] ), .CI(\SUMB[25][29] ), 
        .CO(\CARRYB[26][28] ), .S(\SUMB[26][28] ) );
  FA_X1 S2_26_29 ( .A(\ab[26][29] ), .B(\CARRYB[25][29] ), .CI(\SUMB[25][30] ), 
        .CO(\CARRYB[26][29] ), .S(\SUMB[26][29] ) );
  FA_X1 S3_26_30 ( .A(\ab[26][30] ), .B(\CARRYB[25][30] ), .CI(\ab[25][31] ), 
        .CO(\CARRYB[26][30] ), .S(\SUMB[26][30] ) );
  FA_X1 S1_25_0 ( .A(\ab[25][0] ), .B(\CARRYB[24][0] ), .CI(\SUMB[24][1] ), 
        .CO(\CARRYB[25][0] ), .S(\A1[23] ) );
  FA_X1 S2_25_1 ( .A(\ab[25][1] ), .B(\CARRYB[24][1] ), .CI(\SUMB[24][2] ), 
        .CO(\CARRYB[25][1] ), .S(\SUMB[25][1] ) );
  FA_X1 S2_25_2 ( .A(\ab[25][2] ), .B(\CARRYB[24][2] ), .CI(\SUMB[24][3] ), 
        .CO(\CARRYB[25][2] ), .S(\SUMB[25][2] ) );
  FA_X1 S2_25_3 ( .A(\ab[25][3] ), .B(\CARRYB[24][3] ), .CI(\SUMB[24][4] ), 
        .CO(\CARRYB[25][3] ), .S(\SUMB[25][3] ) );
  FA_X1 S2_25_4 ( .A(\ab[25][4] ), .B(\CARRYB[24][4] ), .CI(\SUMB[24][5] ), 
        .CO(\CARRYB[25][4] ), .S(\SUMB[25][4] ) );
  FA_X1 S2_25_5 ( .A(\ab[25][5] ), .B(\CARRYB[24][5] ), .CI(\SUMB[24][6] ), 
        .CO(\CARRYB[25][5] ), .S(\SUMB[25][5] ) );
  FA_X1 S2_25_6 ( .A(\ab[25][6] ), .B(\CARRYB[24][6] ), .CI(\SUMB[24][7] ), 
        .CO(\CARRYB[25][6] ), .S(\SUMB[25][6] ) );
  FA_X1 S2_25_7 ( .A(\CARRYB[24][7] ), .B(\ab[25][7] ), .CI(\SUMB[24][8] ), 
        .CO(\CARRYB[25][7] ), .S(\SUMB[25][7] ) );
  FA_X1 S2_25_8 ( .A(\CARRYB[24][8] ), .B(\ab[25][8] ), .CI(\SUMB[24][9] ), 
        .CO(\CARRYB[25][8] ), .S(\SUMB[25][8] ) );
  FA_X1 S2_25_11 ( .A(\ab[25][11] ), .B(\CARRYB[24][11] ), .CI(\SUMB[24][12] ), 
        .CO(\CARRYB[25][11] ), .S(\SUMB[25][11] ) );
  FA_X1 S2_25_12 ( .A(\ab[25][12] ), .B(\CARRYB[24][12] ), .CI(\SUMB[24][13] ), 
        .CO(\CARRYB[25][12] ), .S(\SUMB[25][12] ) );
  FA_X1 S2_25_13 ( .A(\ab[25][13] ), .B(\CARRYB[24][13] ), .CI(\SUMB[24][14] ), 
        .CO(\CARRYB[25][13] ), .S(\SUMB[25][13] ) );
  FA_X1 S2_25_14 ( .A(\ab[25][14] ), .B(\CARRYB[24][14] ), .CI(\SUMB[24][15] ), 
        .CO(\CARRYB[25][14] ), .S(\SUMB[25][14] ) );
  FA_X1 S2_25_15 ( .A(\ab[25][15] ), .B(\CARRYB[24][15] ), .CI(\SUMB[24][16] ), 
        .CO(\CARRYB[25][15] ), .S(\SUMB[25][15] ) );
  FA_X1 S2_25_16 ( .A(\ab[25][16] ), .B(\CARRYB[24][16] ), .CI(\SUMB[24][17] ), 
        .CO(\CARRYB[25][16] ), .S(\SUMB[25][16] ) );
  FA_X1 S2_25_17 ( .A(\ab[25][17] ), .B(\CARRYB[24][17] ), .CI(\SUMB[24][18] ), 
        .CO(\CARRYB[25][17] ), .S(\SUMB[25][17] ) );
  FA_X1 S2_25_18 ( .A(\ab[25][18] ), .B(\CARRYB[24][18] ), .CI(\SUMB[24][19] ), 
        .CO(\CARRYB[25][18] ), .S(\SUMB[25][18] ) );
  FA_X1 S2_25_19 ( .A(\ab[25][19] ), .B(\CARRYB[24][19] ), .CI(\SUMB[24][20] ), 
        .CO(\CARRYB[25][19] ), .S(\SUMB[25][19] ) );
  FA_X1 S2_25_20 ( .A(\ab[25][20] ), .B(\CARRYB[24][20] ), .CI(\SUMB[24][21] ), 
        .CO(\CARRYB[25][20] ), .S(\SUMB[25][20] ) );
  FA_X1 S2_25_21 ( .A(\ab[25][21] ), .B(\CARRYB[24][21] ), .CI(\SUMB[24][22] ), 
        .CO(\CARRYB[25][21] ), .S(\SUMB[25][21] ) );
  FA_X1 S2_25_22 ( .A(\ab[25][22] ), .B(\CARRYB[24][22] ), .CI(\SUMB[24][23] ), 
        .CO(\CARRYB[25][22] ), .S(\SUMB[25][22] ) );
  FA_X1 S2_25_23 ( .A(\ab[25][23] ), .B(\CARRYB[24][23] ), .CI(\SUMB[24][24] ), 
        .CO(\CARRYB[25][23] ), .S(\SUMB[25][23] ) );
  FA_X1 S2_25_24 ( .A(\ab[25][24] ), .B(\CARRYB[24][24] ), .CI(\SUMB[24][25] ), 
        .CO(\CARRYB[25][24] ), .S(\SUMB[25][24] ) );
  FA_X1 S2_25_25 ( .A(\ab[25][25] ), .B(\CARRYB[24][25] ), .CI(\SUMB[24][26] ), 
        .CO(\CARRYB[25][25] ), .S(\SUMB[25][25] ) );
  FA_X1 S2_25_26 ( .A(\ab[25][26] ), .B(\CARRYB[24][26] ), .CI(\SUMB[24][27] ), 
        .CO(\CARRYB[25][26] ), .S(\SUMB[25][26] ) );
  FA_X1 S2_25_27 ( .A(\ab[25][27] ), .B(\CARRYB[24][27] ), .CI(\SUMB[24][28] ), 
        .CO(\CARRYB[25][27] ), .S(\SUMB[25][27] ) );
  FA_X1 S2_25_28 ( .A(\ab[25][28] ), .B(\CARRYB[24][28] ), .CI(\SUMB[24][29] ), 
        .CO(\CARRYB[25][28] ), .S(\SUMB[25][28] ) );
  FA_X1 S2_25_29 ( .A(\ab[25][29] ), .B(\CARRYB[24][29] ), .CI(\SUMB[24][30] ), 
        .CO(\CARRYB[25][29] ), .S(\SUMB[25][29] ) );
  FA_X1 S3_25_30 ( .A(\ab[25][30] ), .B(\CARRYB[24][30] ), .CI(\ab[24][31] ), 
        .CO(\CARRYB[25][30] ), .S(\SUMB[25][30] ) );
  FA_X1 S1_24_0 ( .A(\ab[24][0] ), .B(\CARRYB[23][0] ), .CI(\SUMB[23][1] ), 
        .CO(\CARRYB[24][0] ), .S(\A1[22] ) );
  FA_X1 S2_24_1 ( .A(\ab[24][1] ), .B(\CARRYB[23][1] ), .CI(\SUMB[23][2] ), 
        .CO(\CARRYB[24][1] ), .S(\SUMB[24][1] ) );
  FA_X1 S2_24_2 ( .A(\ab[24][2] ), .B(\CARRYB[23][2] ), .CI(\SUMB[23][3] ), 
        .CO(\CARRYB[24][2] ), .S(\SUMB[24][2] ) );
  FA_X1 S2_24_3 ( .A(\ab[24][3] ), .B(\CARRYB[23][3] ), .CI(\SUMB[23][4] ), 
        .CO(\CARRYB[24][3] ), .S(\SUMB[24][3] ) );
  FA_X1 S2_24_4 ( .A(\ab[24][4] ), .B(\CARRYB[23][4] ), .CI(\SUMB[23][5] ), 
        .CO(\CARRYB[24][4] ), .S(\SUMB[24][4] ) );
  FA_X1 S2_24_5 ( .A(\ab[24][5] ), .B(\CARRYB[23][5] ), .CI(\SUMB[23][6] ), 
        .CO(\CARRYB[24][5] ), .S(\SUMB[24][5] ) );
  FA_X1 S2_24_6 ( .A(\ab[24][6] ), .B(\CARRYB[23][6] ), .CI(\SUMB[23][7] ), 
        .CO(\CARRYB[24][6] ), .S(\SUMB[24][6] ) );
  FA_X1 S2_24_7 ( .A(\ab[24][7] ), .B(\CARRYB[23][7] ), .CI(\SUMB[23][8] ), 
        .CO(\CARRYB[24][7] ), .S(\SUMB[24][7] ) );
  FA_X1 S2_24_8 ( .A(\ab[24][8] ), .B(\CARRYB[23][8] ), .CI(\SUMB[23][9] ), 
        .CO(\CARRYB[24][8] ), .S(\SUMB[24][8] ) );
  FA_X1 S2_24_9 ( .A(\CARRYB[23][9] ), .B(\ab[24][9] ), .CI(\SUMB[23][10] ), 
        .CO(\CARRYB[24][9] ), .S(\SUMB[24][9] ) );
  FA_X1 S2_24_12 ( .A(\ab[24][12] ), .B(\CARRYB[23][12] ), .CI(\SUMB[23][13] ), 
        .CO(\CARRYB[24][12] ), .S(\SUMB[24][12] ) );
  FA_X1 S2_24_13 ( .A(\ab[24][13] ), .B(\CARRYB[23][13] ), .CI(\SUMB[23][14] ), 
        .CO(\CARRYB[24][13] ), .S(\SUMB[24][13] ) );
  FA_X1 S2_24_14 ( .A(\ab[24][14] ), .B(\CARRYB[23][14] ), .CI(\SUMB[23][15] ), 
        .CO(\CARRYB[24][14] ), .S(\SUMB[24][14] ) );
  FA_X1 S2_24_15 ( .A(\ab[24][15] ), .B(\CARRYB[23][15] ), .CI(\SUMB[23][16] ), 
        .CO(\CARRYB[24][15] ), .S(\SUMB[24][15] ) );
  FA_X1 S2_24_16 ( .A(\ab[24][16] ), .B(\CARRYB[23][16] ), .CI(\SUMB[23][17] ), 
        .CO(\CARRYB[24][16] ), .S(\SUMB[24][16] ) );
  FA_X1 S2_24_17 ( .A(\ab[24][17] ), .B(\CARRYB[23][17] ), .CI(\SUMB[23][18] ), 
        .CO(\CARRYB[24][17] ), .S(\SUMB[24][17] ) );
  FA_X1 S2_24_18 ( .A(\ab[24][18] ), .B(\CARRYB[23][18] ), .CI(\SUMB[23][19] ), 
        .CO(\CARRYB[24][18] ), .S(\SUMB[24][18] ) );
  FA_X1 S2_24_19 ( .A(\ab[24][19] ), .B(\CARRYB[23][19] ), .CI(\SUMB[23][20] ), 
        .CO(\CARRYB[24][19] ), .S(\SUMB[24][19] ) );
  FA_X1 S2_24_20 ( .A(\ab[24][20] ), .B(\CARRYB[23][20] ), .CI(\SUMB[23][21] ), 
        .CO(\CARRYB[24][20] ), .S(\SUMB[24][20] ) );
  FA_X1 S2_24_21 ( .A(\ab[24][21] ), .B(\CARRYB[23][21] ), .CI(\SUMB[23][22] ), 
        .CO(\CARRYB[24][21] ), .S(\SUMB[24][21] ) );
  FA_X1 S2_24_22 ( .A(\ab[24][22] ), .B(\CARRYB[23][22] ), .CI(\SUMB[23][23] ), 
        .CO(\CARRYB[24][22] ), .S(\SUMB[24][22] ) );
  FA_X1 S2_24_23 ( .A(\ab[24][23] ), .B(\CARRYB[23][23] ), .CI(\SUMB[23][24] ), 
        .CO(\CARRYB[24][23] ), .S(\SUMB[24][23] ) );
  FA_X1 S2_24_24 ( .A(\ab[24][24] ), .B(\CARRYB[23][24] ), .CI(\SUMB[23][25] ), 
        .CO(\CARRYB[24][24] ), .S(\SUMB[24][24] ) );
  FA_X1 S2_24_25 ( .A(\ab[24][25] ), .B(\CARRYB[23][25] ), .CI(\SUMB[23][26] ), 
        .CO(\CARRYB[24][25] ), .S(\SUMB[24][25] ) );
  FA_X1 S2_24_26 ( .A(\ab[24][26] ), .B(\CARRYB[23][26] ), .CI(\SUMB[23][27] ), 
        .CO(\CARRYB[24][26] ), .S(\SUMB[24][26] ) );
  FA_X1 S2_24_27 ( .A(\ab[24][27] ), .B(\CARRYB[23][27] ), .CI(\SUMB[23][28] ), 
        .CO(\CARRYB[24][27] ), .S(\SUMB[24][27] ) );
  FA_X1 S2_24_28 ( .A(\ab[24][28] ), .B(\CARRYB[23][28] ), .CI(\SUMB[23][29] ), 
        .CO(\CARRYB[24][28] ), .S(\SUMB[24][28] ) );
  FA_X1 S2_24_29 ( .A(\ab[24][29] ), .B(\CARRYB[23][29] ), .CI(\SUMB[23][30] ), 
        .CO(\CARRYB[24][29] ), .S(\SUMB[24][29] ) );
  FA_X1 S3_24_30 ( .A(\ab[24][30] ), .B(\CARRYB[23][30] ), .CI(\ab[23][31] ), 
        .CO(\CARRYB[24][30] ), .S(\SUMB[24][30] ) );
  FA_X1 S1_23_0 ( .A(\ab[23][0] ), .B(\CARRYB[22][0] ), .CI(\SUMB[22][1] ), 
        .CO(\CARRYB[23][0] ), .S(\A1[21] ) );
  FA_X1 S2_23_1 ( .A(\ab[23][1] ), .B(\CARRYB[22][1] ), .CI(\SUMB[22][2] ), 
        .CO(\CARRYB[23][1] ), .S(\SUMB[23][1] ) );
  FA_X1 S2_23_2 ( .A(\ab[23][2] ), .B(\CARRYB[22][2] ), .CI(\SUMB[22][3] ), 
        .CO(\CARRYB[23][2] ), .S(\SUMB[23][2] ) );
  FA_X1 S2_23_3 ( .A(\ab[23][3] ), .B(\CARRYB[22][3] ), .CI(\SUMB[22][4] ), 
        .CO(\CARRYB[23][3] ), .S(\SUMB[23][3] ) );
  FA_X1 S2_23_4 ( .A(\ab[23][4] ), .B(\CARRYB[22][4] ), .CI(\SUMB[22][5] ), 
        .CO(\CARRYB[23][4] ), .S(\SUMB[23][4] ) );
  FA_X1 S2_23_5 ( .A(\ab[23][5] ), .B(\CARRYB[22][5] ), .CI(\SUMB[22][6] ), 
        .CO(\CARRYB[23][5] ), .S(\SUMB[23][5] ) );
  FA_X1 S2_23_6 ( .A(\ab[23][6] ), .B(\CARRYB[22][6] ), .CI(\SUMB[22][7] ), 
        .CO(\CARRYB[23][6] ), .S(\SUMB[23][6] ) );
  FA_X1 S2_23_7 ( .A(\ab[23][7] ), .B(\CARRYB[22][7] ), .CI(\SUMB[22][8] ), 
        .CO(\CARRYB[23][7] ), .S(\SUMB[23][7] ) );
  FA_X1 S2_23_8 ( .A(\ab[23][8] ), .B(\CARRYB[22][8] ), .CI(\SUMB[22][9] ), 
        .CO(\CARRYB[23][8] ), .S(\SUMB[23][8] ) );
  FA_X1 S2_23_9 ( .A(\CARRYB[22][9] ), .B(\ab[23][9] ), .CI(\SUMB[22][10] ), 
        .CO(\CARRYB[23][9] ), .S(\SUMB[23][9] ) );
  FA_X1 S2_23_10 ( .A(\ab[23][10] ), .B(\CARRYB[22][10] ), .CI(\SUMB[22][11] ), 
        .CO(\CARRYB[23][10] ), .S(\SUMB[23][10] ) );
  FA_X1 S2_23_13 ( .A(\ab[23][13] ), .B(\CARRYB[22][13] ), .CI(\SUMB[22][14] ), 
        .CO(\CARRYB[23][13] ), .S(\SUMB[23][13] ) );
  FA_X1 S2_23_14 ( .A(\ab[23][14] ), .B(\CARRYB[22][14] ), .CI(\SUMB[22][15] ), 
        .CO(\CARRYB[23][14] ), .S(\SUMB[23][14] ) );
  FA_X1 S2_23_15 ( .A(\ab[23][15] ), .B(\CARRYB[22][15] ), .CI(\SUMB[22][16] ), 
        .CO(\CARRYB[23][15] ), .S(\SUMB[23][15] ) );
  FA_X1 S2_23_16 ( .A(\ab[23][16] ), .B(\CARRYB[22][16] ), .CI(\SUMB[22][17] ), 
        .CO(\CARRYB[23][16] ), .S(\SUMB[23][16] ) );
  FA_X1 S2_23_17 ( .A(\ab[23][17] ), .B(\CARRYB[22][17] ), .CI(\SUMB[22][18] ), 
        .CO(\CARRYB[23][17] ), .S(\SUMB[23][17] ) );
  FA_X1 S2_23_18 ( .A(\ab[23][18] ), .B(\CARRYB[22][18] ), .CI(\SUMB[22][19] ), 
        .CO(\CARRYB[23][18] ), .S(\SUMB[23][18] ) );
  FA_X1 S2_23_19 ( .A(\ab[23][19] ), .B(\CARRYB[22][19] ), .CI(\SUMB[22][20] ), 
        .CO(\CARRYB[23][19] ), .S(\SUMB[23][19] ) );
  FA_X1 S2_23_20 ( .A(\ab[23][20] ), .B(\CARRYB[22][20] ), .CI(\SUMB[22][21] ), 
        .CO(\CARRYB[23][20] ), .S(\SUMB[23][20] ) );
  FA_X1 S2_23_21 ( .A(\ab[23][21] ), .B(\CARRYB[22][21] ), .CI(\SUMB[22][22] ), 
        .CO(\CARRYB[23][21] ), .S(\SUMB[23][21] ) );
  FA_X1 S2_23_22 ( .A(\ab[23][22] ), .B(\CARRYB[22][22] ), .CI(\SUMB[22][23] ), 
        .CO(\CARRYB[23][22] ), .S(\SUMB[23][22] ) );
  FA_X1 S2_23_23 ( .A(\ab[23][23] ), .B(\CARRYB[22][23] ), .CI(\SUMB[22][24] ), 
        .CO(\CARRYB[23][23] ), .S(\SUMB[23][23] ) );
  FA_X1 S2_23_24 ( .A(\ab[23][24] ), .B(\CARRYB[22][24] ), .CI(\SUMB[22][25] ), 
        .CO(\CARRYB[23][24] ), .S(\SUMB[23][24] ) );
  FA_X1 S2_23_25 ( .A(\ab[23][25] ), .B(\CARRYB[22][25] ), .CI(\SUMB[22][26] ), 
        .CO(\CARRYB[23][25] ), .S(\SUMB[23][25] ) );
  FA_X1 S2_23_26 ( .A(\ab[23][26] ), .B(\CARRYB[22][26] ), .CI(\SUMB[22][27] ), 
        .CO(\CARRYB[23][26] ), .S(\SUMB[23][26] ) );
  FA_X1 S2_23_27 ( .A(\ab[23][27] ), .B(\CARRYB[22][27] ), .CI(\SUMB[22][28] ), 
        .CO(\CARRYB[23][27] ), .S(\SUMB[23][27] ) );
  FA_X1 S2_23_28 ( .A(\ab[23][28] ), .B(\CARRYB[22][28] ), .CI(\SUMB[22][29] ), 
        .CO(\CARRYB[23][28] ), .S(\SUMB[23][28] ) );
  FA_X1 S2_23_29 ( .A(\ab[23][29] ), .B(\CARRYB[22][29] ), .CI(\SUMB[22][30] ), 
        .CO(\CARRYB[23][29] ), .S(\SUMB[23][29] ) );
  FA_X1 S3_23_30 ( .A(\ab[23][30] ), .B(\CARRYB[22][30] ), .CI(\ab[22][31] ), 
        .CO(\CARRYB[23][30] ), .S(\SUMB[23][30] ) );
  FA_X1 S1_22_0 ( .A(\ab[22][0] ), .B(\CARRYB[21][0] ), .CI(\SUMB[21][1] ), 
        .CO(\CARRYB[22][0] ), .S(\A1[20] ) );
  FA_X1 S2_22_1 ( .A(\ab[22][1] ), .B(\CARRYB[21][1] ), .CI(\SUMB[21][2] ), 
        .CO(\CARRYB[22][1] ), .S(\SUMB[22][1] ) );
  FA_X1 S2_22_2 ( .A(\ab[22][2] ), .B(\CARRYB[21][2] ), .CI(\SUMB[21][3] ), 
        .CO(\CARRYB[22][2] ), .S(\SUMB[22][2] ) );
  FA_X1 S2_22_3 ( .A(\ab[22][3] ), .B(\CARRYB[21][3] ), .CI(\SUMB[21][4] ), 
        .CO(\CARRYB[22][3] ), .S(\SUMB[22][3] ) );
  FA_X1 S2_22_4 ( .A(\ab[22][4] ), .B(\CARRYB[21][4] ), .CI(\SUMB[21][5] ), 
        .CO(\CARRYB[22][4] ), .S(\SUMB[22][4] ) );
  FA_X1 S2_22_5 ( .A(\ab[22][5] ), .B(\CARRYB[21][5] ), .CI(\SUMB[21][6] ), 
        .CO(\CARRYB[22][5] ), .S(\SUMB[22][5] ) );
  FA_X1 S2_22_6 ( .A(\ab[22][6] ), .B(\CARRYB[21][6] ), .CI(\SUMB[21][7] ), 
        .CO(\CARRYB[22][6] ), .S(\SUMB[22][6] ) );
  FA_X1 S2_22_7 ( .A(\ab[22][7] ), .B(\CARRYB[21][7] ), .CI(\SUMB[21][8] ), 
        .CO(\CARRYB[22][7] ), .S(\SUMB[22][7] ) );
  FA_X1 S2_22_8 ( .A(\ab[22][8] ), .B(\CARRYB[21][8] ), .CI(\SUMB[21][9] ), 
        .CO(\CARRYB[22][8] ), .S(\SUMB[22][8] ) );
  FA_X1 S2_22_9 ( .A(\ab[22][9] ), .B(\CARRYB[21][9] ), .CI(\SUMB[21][10] ), 
        .CO(\CARRYB[22][9] ), .S(\SUMB[22][9] ) );
  FA_X1 S2_22_10 ( .A(\ab[22][10] ), .B(\CARRYB[21][10] ), .CI(\SUMB[21][11] ), 
        .CO(\CARRYB[22][10] ), .S(\SUMB[22][10] ) );
  FA_X1 S2_22_11 ( .A(\CARRYB[21][11] ), .B(\ab[22][11] ), .CI(\SUMB[21][12] ), 
        .CO(\CARRYB[22][11] ), .S(\SUMB[22][11] ) );
  FA_X1 S2_22_14 ( .A(\ab[22][14] ), .B(\CARRYB[21][14] ), .CI(\SUMB[21][15] ), 
        .CO(\CARRYB[22][14] ), .S(\SUMB[22][14] ) );
  FA_X1 S2_22_15 ( .A(\ab[22][15] ), .B(\CARRYB[21][15] ), .CI(\SUMB[21][16] ), 
        .CO(\CARRYB[22][15] ), .S(\SUMB[22][15] ) );
  FA_X1 S2_22_16 ( .A(\ab[22][16] ), .B(\CARRYB[21][16] ), .CI(\SUMB[21][17] ), 
        .CO(\CARRYB[22][16] ), .S(\SUMB[22][16] ) );
  FA_X1 S2_22_17 ( .A(\ab[22][17] ), .B(\CARRYB[21][17] ), .CI(\SUMB[21][18] ), 
        .CO(\CARRYB[22][17] ), .S(\SUMB[22][17] ) );
  FA_X1 S2_22_18 ( .A(\ab[22][18] ), .B(\CARRYB[21][18] ), .CI(\SUMB[21][19] ), 
        .CO(\CARRYB[22][18] ), .S(\SUMB[22][18] ) );
  FA_X1 S2_22_19 ( .A(\ab[22][19] ), .B(\CARRYB[21][19] ), .CI(\SUMB[21][20] ), 
        .CO(\CARRYB[22][19] ), .S(\SUMB[22][19] ) );
  FA_X1 S2_22_20 ( .A(\ab[22][20] ), .B(\CARRYB[21][20] ), .CI(\SUMB[21][21] ), 
        .CO(\CARRYB[22][20] ), .S(\SUMB[22][20] ) );
  FA_X1 S2_22_21 ( .A(\ab[22][21] ), .B(\CARRYB[21][21] ), .CI(\SUMB[21][22] ), 
        .CO(\CARRYB[22][21] ), .S(\SUMB[22][21] ) );
  FA_X1 S2_22_22 ( .A(\ab[22][22] ), .B(\CARRYB[21][22] ), .CI(\SUMB[21][23] ), 
        .CO(\CARRYB[22][22] ), .S(\SUMB[22][22] ) );
  FA_X1 S2_22_23 ( .A(\ab[22][23] ), .B(\CARRYB[21][23] ), .CI(\SUMB[21][24] ), 
        .CO(\CARRYB[22][23] ), .S(\SUMB[22][23] ) );
  FA_X1 S2_22_24 ( .A(\ab[22][24] ), .B(\CARRYB[21][24] ), .CI(\SUMB[21][25] ), 
        .CO(\CARRYB[22][24] ), .S(\SUMB[22][24] ) );
  FA_X1 S2_22_25 ( .A(\ab[22][25] ), .B(\CARRYB[21][25] ), .CI(\SUMB[21][26] ), 
        .CO(\CARRYB[22][25] ), .S(\SUMB[22][25] ) );
  FA_X1 S2_22_26 ( .A(\ab[22][26] ), .B(\CARRYB[21][26] ), .CI(\SUMB[21][27] ), 
        .CO(\CARRYB[22][26] ), .S(\SUMB[22][26] ) );
  FA_X1 S2_22_27 ( .A(\ab[22][27] ), .B(\CARRYB[21][27] ), .CI(\SUMB[21][28] ), 
        .CO(\CARRYB[22][27] ), .S(\SUMB[22][27] ) );
  FA_X1 S2_22_28 ( .A(\ab[22][28] ), .B(\CARRYB[21][28] ), .CI(\SUMB[21][29] ), 
        .CO(\CARRYB[22][28] ), .S(\SUMB[22][28] ) );
  FA_X1 S2_22_29 ( .A(\ab[22][29] ), .B(\CARRYB[21][29] ), .CI(\SUMB[21][30] ), 
        .CO(\CARRYB[22][29] ), .S(\SUMB[22][29] ) );
  FA_X1 S3_22_30 ( .A(\ab[22][30] ), .B(\CARRYB[21][30] ), .CI(\ab[21][31] ), 
        .CO(\CARRYB[22][30] ), .S(\SUMB[22][30] ) );
  FA_X1 S1_21_0 ( .A(\ab[21][0] ), .B(\CARRYB[20][0] ), .CI(\SUMB[20][1] ), 
        .CO(\CARRYB[21][0] ), .S(\A1[19] ) );
  FA_X1 S2_21_1 ( .A(\ab[21][1] ), .B(\CARRYB[20][1] ), .CI(\SUMB[20][2] ), 
        .CO(\CARRYB[21][1] ), .S(\SUMB[21][1] ) );
  FA_X1 S2_21_2 ( .A(\ab[21][2] ), .B(\CARRYB[20][2] ), .CI(\SUMB[20][3] ), 
        .CO(\CARRYB[21][2] ), .S(\SUMB[21][2] ) );
  FA_X1 S2_21_3 ( .A(\ab[21][3] ), .B(\CARRYB[20][3] ), .CI(\SUMB[20][4] ), 
        .CO(\CARRYB[21][3] ), .S(\SUMB[21][3] ) );
  FA_X1 S2_21_4 ( .A(\ab[21][4] ), .B(\CARRYB[20][4] ), .CI(\SUMB[20][5] ), 
        .CO(\CARRYB[21][4] ), .S(\SUMB[21][4] ) );
  FA_X1 S2_21_5 ( .A(\ab[21][5] ), .B(\CARRYB[20][5] ), .CI(\SUMB[20][6] ), 
        .CO(\CARRYB[21][5] ), .S(\SUMB[21][5] ) );
  FA_X1 S2_21_6 ( .A(\ab[21][6] ), .B(\CARRYB[20][6] ), .CI(\SUMB[20][7] ), 
        .CO(\CARRYB[21][6] ), .S(\SUMB[21][6] ) );
  FA_X1 S2_21_7 ( .A(\ab[21][7] ), .B(\CARRYB[20][7] ), .CI(\SUMB[20][8] ), 
        .CO(\CARRYB[21][7] ), .S(\SUMB[21][7] ) );
  FA_X1 S2_21_8 ( .A(\ab[21][8] ), .B(\CARRYB[20][8] ), .CI(\SUMB[20][9] ), 
        .CO(\CARRYB[21][8] ), .S(\SUMB[21][8] ) );
  FA_X1 S2_21_9 ( .A(\ab[21][9] ), .B(\CARRYB[20][9] ), .CI(\SUMB[20][10] ), 
        .CO(\CARRYB[21][9] ), .S(\SUMB[21][9] ) );
  FA_X1 S2_21_10 ( .A(\ab[21][10] ), .B(\CARRYB[20][10] ), .CI(\SUMB[20][11] ), 
        .CO(\CARRYB[21][10] ), .S(\SUMB[21][10] ) );
  FA_X1 S2_21_11 ( .A(\CARRYB[20][11] ), .B(\ab[21][11] ), .CI(\SUMB[20][12] ), 
        .CO(\CARRYB[21][11] ), .S(\SUMB[21][11] ) );
  FA_X1 S2_21_12 ( .A(\ab[21][12] ), .B(\CARRYB[20][12] ), .CI(\SUMB[20][13] ), 
        .CO(\CARRYB[21][12] ), .S(\SUMB[21][12] ) );
  FA_X1 S2_21_15 ( .A(\ab[21][15] ), .B(\CARRYB[20][15] ), .CI(\SUMB[20][16] ), 
        .CO(\CARRYB[21][15] ), .S(\SUMB[21][15] ) );
  FA_X1 S2_21_16 ( .A(\ab[21][16] ), .B(\CARRYB[20][16] ), .CI(\SUMB[20][17] ), 
        .CO(\CARRYB[21][16] ), .S(\SUMB[21][16] ) );
  FA_X1 S2_21_17 ( .A(\ab[21][17] ), .B(\CARRYB[20][17] ), .CI(\SUMB[20][18] ), 
        .CO(\CARRYB[21][17] ), .S(\SUMB[21][17] ) );
  FA_X1 S2_21_18 ( .A(\ab[21][18] ), .B(\CARRYB[20][18] ), .CI(\SUMB[20][19] ), 
        .CO(\CARRYB[21][18] ), .S(\SUMB[21][18] ) );
  FA_X1 S2_21_19 ( .A(\ab[21][19] ), .B(\CARRYB[20][19] ), .CI(\SUMB[20][20] ), 
        .CO(\CARRYB[21][19] ), .S(\SUMB[21][19] ) );
  FA_X1 S2_21_20 ( .A(\ab[21][20] ), .B(\CARRYB[20][20] ), .CI(\SUMB[20][21] ), 
        .CO(\CARRYB[21][20] ), .S(\SUMB[21][20] ) );
  FA_X1 S2_21_21 ( .A(\ab[21][21] ), .B(\CARRYB[20][21] ), .CI(\SUMB[20][22] ), 
        .CO(\CARRYB[21][21] ), .S(\SUMB[21][21] ) );
  FA_X1 S2_21_22 ( .A(\ab[21][22] ), .B(\CARRYB[20][22] ), .CI(\SUMB[20][23] ), 
        .CO(\CARRYB[21][22] ), .S(\SUMB[21][22] ) );
  FA_X1 S2_21_23 ( .A(\ab[21][23] ), .B(\CARRYB[20][23] ), .CI(\SUMB[20][24] ), 
        .CO(\CARRYB[21][23] ), .S(\SUMB[21][23] ) );
  FA_X1 S2_21_24 ( .A(\ab[21][24] ), .B(\CARRYB[20][24] ), .CI(\SUMB[20][25] ), 
        .CO(\CARRYB[21][24] ), .S(\SUMB[21][24] ) );
  FA_X1 S2_21_25 ( .A(\ab[21][25] ), .B(\CARRYB[20][25] ), .CI(\SUMB[20][26] ), 
        .CO(\CARRYB[21][25] ), .S(\SUMB[21][25] ) );
  FA_X1 S2_21_26 ( .A(\ab[21][26] ), .B(\CARRYB[20][26] ), .CI(\SUMB[20][27] ), 
        .CO(\CARRYB[21][26] ), .S(\SUMB[21][26] ) );
  FA_X1 S2_21_27 ( .A(\ab[21][27] ), .B(\CARRYB[20][27] ), .CI(\SUMB[20][28] ), 
        .CO(\CARRYB[21][27] ), .S(\SUMB[21][27] ) );
  FA_X1 S2_21_28 ( .A(\ab[21][28] ), .B(\CARRYB[20][28] ), .CI(\SUMB[20][29] ), 
        .CO(\CARRYB[21][28] ), .S(\SUMB[21][28] ) );
  FA_X1 S2_21_29 ( .A(\ab[21][29] ), .B(\CARRYB[20][29] ), .CI(\SUMB[20][30] ), 
        .CO(\CARRYB[21][29] ), .S(\SUMB[21][29] ) );
  FA_X1 S3_21_30 ( .A(\ab[21][30] ), .B(\CARRYB[20][30] ), .CI(\ab[20][31] ), 
        .CO(\CARRYB[21][30] ), .S(\SUMB[21][30] ) );
  FA_X1 S1_20_0 ( .A(\ab[20][0] ), .B(\CARRYB[19][0] ), .CI(\SUMB[19][1] ), 
        .CO(\CARRYB[20][0] ), .S(\A1[18] ) );
  FA_X1 S2_20_1 ( .A(\ab[20][1] ), .B(\CARRYB[19][1] ), .CI(\SUMB[19][2] ), 
        .CO(\CARRYB[20][1] ), .S(\SUMB[20][1] ) );
  FA_X1 S2_20_2 ( .A(\ab[20][2] ), .B(\CARRYB[19][2] ), .CI(\SUMB[19][3] ), 
        .CO(\CARRYB[20][2] ), .S(\SUMB[20][2] ) );
  FA_X1 S2_20_3 ( .A(\ab[20][3] ), .B(\CARRYB[19][3] ), .CI(\SUMB[19][4] ), 
        .CO(\CARRYB[20][3] ), .S(\SUMB[20][3] ) );
  FA_X1 S2_20_4 ( .A(\ab[20][4] ), .B(\CARRYB[19][4] ), .CI(\SUMB[19][5] ), 
        .CO(\CARRYB[20][4] ), .S(\SUMB[20][4] ) );
  FA_X1 S2_20_5 ( .A(\ab[20][5] ), .B(\CARRYB[19][5] ), .CI(\SUMB[19][6] ), 
        .CO(\CARRYB[20][5] ), .S(\SUMB[20][5] ) );
  FA_X1 S2_20_6 ( .A(\ab[20][6] ), .B(\CARRYB[19][6] ), .CI(\SUMB[19][7] ), 
        .CO(\CARRYB[20][6] ), .S(\SUMB[20][6] ) );
  FA_X1 S2_20_7 ( .A(\ab[20][7] ), .B(\CARRYB[19][7] ), .CI(\SUMB[19][8] ), 
        .CO(\CARRYB[20][7] ), .S(\SUMB[20][7] ) );
  FA_X1 S2_20_8 ( .A(\ab[20][8] ), .B(\CARRYB[19][8] ), .CI(\SUMB[19][9] ), 
        .CO(\CARRYB[20][8] ), .S(\SUMB[20][8] ) );
  FA_X1 S2_20_9 ( .A(\ab[20][9] ), .B(\CARRYB[19][9] ), .CI(\SUMB[19][10] ), 
        .CO(\CARRYB[20][9] ), .S(\SUMB[20][9] ) );
  FA_X1 S2_20_10 ( .A(\ab[20][10] ), .B(\CARRYB[19][10] ), .CI(\SUMB[19][11] ), 
        .CO(\CARRYB[20][10] ), .S(\SUMB[20][10] ) );
  FA_X1 S2_20_11 ( .A(\ab[20][11] ), .B(\CARRYB[19][11] ), .CI(\SUMB[19][12] ), 
        .CO(\CARRYB[20][11] ), .S(\SUMB[20][11] ) );
  FA_X1 S2_20_12 ( .A(\ab[20][12] ), .B(\CARRYB[19][12] ), .CI(\SUMB[19][13] ), 
        .CO(\CARRYB[20][12] ), .S(\SUMB[20][12] ) );
  FA_X1 S2_20_13 ( .A(\CARRYB[19][13] ), .B(\ab[20][13] ), .CI(\SUMB[19][14] ), 
        .CO(\CARRYB[20][13] ), .S(\SUMB[20][13] ) );
  FA_X1 S2_20_16 ( .A(\ab[20][16] ), .B(\CARRYB[19][16] ), .CI(\SUMB[19][17] ), 
        .CO(\CARRYB[20][16] ), .S(\SUMB[20][16] ) );
  FA_X1 S2_20_17 ( .A(\ab[20][17] ), .B(\CARRYB[19][17] ), .CI(\SUMB[19][18] ), 
        .CO(\CARRYB[20][17] ), .S(\SUMB[20][17] ) );
  FA_X1 S2_20_18 ( .A(\ab[20][18] ), .B(\CARRYB[19][18] ), .CI(\SUMB[19][19] ), 
        .CO(\CARRYB[20][18] ), .S(\SUMB[20][18] ) );
  FA_X1 S2_20_19 ( .A(\ab[20][19] ), .B(\CARRYB[19][19] ), .CI(\SUMB[19][20] ), 
        .CO(\CARRYB[20][19] ), .S(\SUMB[20][19] ) );
  FA_X1 S2_20_20 ( .A(\ab[20][20] ), .B(\CARRYB[19][20] ), .CI(\SUMB[19][21] ), 
        .CO(\CARRYB[20][20] ), .S(\SUMB[20][20] ) );
  FA_X1 S2_20_21 ( .A(\ab[20][21] ), .B(\CARRYB[19][21] ), .CI(\SUMB[19][22] ), 
        .CO(\CARRYB[20][21] ), .S(\SUMB[20][21] ) );
  FA_X1 S2_20_22 ( .A(\ab[20][22] ), .B(\CARRYB[19][22] ), .CI(\SUMB[19][23] ), 
        .CO(\CARRYB[20][22] ), .S(\SUMB[20][22] ) );
  FA_X1 S2_20_23 ( .A(\ab[20][23] ), .B(\CARRYB[19][23] ), .CI(\SUMB[19][24] ), 
        .CO(\CARRYB[20][23] ), .S(\SUMB[20][23] ) );
  FA_X1 S2_20_24 ( .A(\ab[20][24] ), .B(\CARRYB[19][24] ), .CI(\SUMB[19][25] ), 
        .CO(\CARRYB[20][24] ), .S(\SUMB[20][24] ) );
  FA_X1 S2_20_25 ( .A(\ab[20][25] ), .B(\CARRYB[19][25] ), .CI(\SUMB[19][26] ), 
        .CO(\CARRYB[20][25] ), .S(\SUMB[20][25] ) );
  FA_X1 S2_20_26 ( .A(\ab[20][26] ), .B(\CARRYB[19][26] ), .CI(\SUMB[19][27] ), 
        .CO(\CARRYB[20][26] ), .S(\SUMB[20][26] ) );
  FA_X1 S2_20_27 ( .A(\ab[20][27] ), .B(\CARRYB[19][27] ), .CI(\SUMB[19][28] ), 
        .CO(\CARRYB[20][27] ), .S(\SUMB[20][27] ) );
  FA_X1 S2_20_28 ( .A(\ab[20][28] ), .B(\CARRYB[19][28] ), .CI(\SUMB[19][29] ), 
        .CO(\CARRYB[20][28] ), .S(\SUMB[20][28] ) );
  FA_X1 S2_20_29 ( .A(\ab[20][29] ), .B(\CARRYB[19][29] ), .CI(\SUMB[19][30] ), 
        .CO(\CARRYB[20][29] ), .S(\SUMB[20][29] ) );
  FA_X1 S3_20_30 ( .A(\ab[20][30] ), .B(\CARRYB[19][30] ), .CI(\ab[19][31] ), 
        .CO(\CARRYB[20][30] ), .S(\SUMB[20][30] ) );
  FA_X1 S1_19_0 ( .A(\ab[19][0] ), .B(\CARRYB[18][0] ), .CI(\SUMB[18][1] ), 
        .CO(\CARRYB[19][0] ), .S(\A1[17] ) );
  FA_X1 S2_19_1 ( .A(\ab[19][1] ), .B(\CARRYB[18][1] ), .CI(\SUMB[18][2] ), 
        .CO(\CARRYB[19][1] ), .S(\SUMB[19][1] ) );
  FA_X1 S2_19_2 ( .A(\ab[19][2] ), .B(\CARRYB[18][2] ), .CI(\SUMB[18][3] ), 
        .CO(\CARRYB[19][2] ), .S(\SUMB[19][2] ) );
  FA_X1 S2_19_3 ( .A(\ab[19][3] ), .B(\CARRYB[18][3] ), .CI(\SUMB[18][4] ), 
        .CO(\CARRYB[19][3] ), .S(\SUMB[19][3] ) );
  FA_X1 S2_19_4 ( .A(\ab[19][4] ), .B(\CARRYB[18][4] ), .CI(\SUMB[18][5] ), 
        .CO(\CARRYB[19][4] ), .S(\SUMB[19][4] ) );
  FA_X1 S2_19_5 ( .A(\ab[19][5] ), .B(\CARRYB[18][5] ), .CI(\SUMB[18][6] ), 
        .CO(\CARRYB[19][5] ), .S(\SUMB[19][5] ) );
  FA_X1 S2_19_6 ( .A(\ab[19][6] ), .B(\CARRYB[18][6] ), .CI(\SUMB[18][7] ), 
        .CO(\CARRYB[19][6] ), .S(\SUMB[19][6] ) );
  FA_X1 S2_19_7 ( .A(\ab[19][7] ), .B(\CARRYB[18][7] ), .CI(\SUMB[18][8] ), 
        .CO(\CARRYB[19][7] ), .S(\SUMB[19][7] ) );
  FA_X1 S2_19_8 ( .A(\ab[19][8] ), .B(\CARRYB[18][8] ), .CI(\SUMB[18][9] ), 
        .CO(\CARRYB[19][8] ), .S(\SUMB[19][8] ) );
  FA_X1 S2_19_9 ( .A(\ab[19][9] ), .B(\CARRYB[18][9] ), .CI(\SUMB[18][10] ), 
        .CO(\CARRYB[19][9] ), .S(\SUMB[19][9] ) );
  FA_X1 S2_19_10 ( .A(\ab[19][10] ), .B(\CARRYB[18][10] ), .CI(\SUMB[18][11] ), 
        .CO(\CARRYB[19][10] ), .S(\SUMB[19][10] ) );
  FA_X1 S2_19_11 ( .A(\ab[19][11] ), .B(\CARRYB[18][11] ), .CI(\SUMB[18][12] ), 
        .CO(\CARRYB[19][11] ), .S(\SUMB[19][11] ) );
  FA_X1 S2_19_12 ( .A(\ab[19][12] ), .B(\CARRYB[18][12] ), .CI(\SUMB[18][13] ), 
        .CO(\CARRYB[19][12] ), .S(\SUMB[19][12] ) );
  FA_X1 S2_19_13 ( .A(\CARRYB[18][13] ), .B(\ab[19][13] ), .CI(\SUMB[18][14] ), 
        .CO(\CARRYB[19][13] ), .S(\SUMB[19][13] ) );
  FA_X1 S2_19_17 ( .A(\ab[19][17] ), .B(\CARRYB[18][17] ), .CI(\SUMB[18][18] ), 
        .CO(\CARRYB[19][17] ), .S(\SUMB[19][17] ) );
  FA_X1 S2_19_18 ( .A(\ab[19][18] ), .B(\CARRYB[18][18] ), .CI(\SUMB[18][19] ), 
        .CO(\CARRYB[19][18] ), .S(\SUMB[19][18] ) );
  FA_X1 S2_19_19 ( .A(\ab[19][19] ), .B(\CARRYB[18][19] ), .CI(\SUMB[18][20] ), 
        .CO(\CARRYB[19][19] ), .S(\SUMB[19][19] ) );
  FA_X1 S2_19_20 ( .A(\ab[19][20] ), .B(\CARRYB[18][20] ), .CI(\SUMB[18][21] ), 
        .CO(\CARRYB[19][20] ), .S(\SUMB[19][20] ) );
  FA_X1 S2_19_21 ( .A(\ab[19][21] ), .B(\CARRYB[18][21] ), .CI(\SUMB[18][22] ), 
        .CO(\CARRYB[19][21] ), .S(\SUMB[19][21] ) );
  FA_X1 S2_19_22 ( .A(\ab[19][22] ), .B(\CARRYB[18][22] ), .CI(\SUMB[18][23] ), 
        .CO(\CARRYB[19][22] ), .S(\SUMB[19][22] ) );
  FA_X1 S2_19_23 ( .A(\ab[19][23] ), .B(\CARRYB[18][23] ), .CI(\SUMB[18][24] ), 
        .CO(\CARRYB[19][23] ), .S(\SUMB[19][23] ) );
  FA_X1 S2_19_24 ( .A(\ab[19][24] ), .B(\CARRYB[18][24] ), .CI(\SUMB[18][25] ), 
        .CO(\CARRYB[19][24] ), .S(\SUMB[19][24] ) );
  FA_X1 S2_19_25 ( .A(\ab[19][25] ), .B(\CARRYB[18][25] ), .CI(\SUMB[18][26] ), 
        .CO(\CARRYB[19][25] ), .S(\SUMB[19][25] ) );
  FA_X1 S2_19_26 ( .A(\ab[19][26] ), .B(\CARRYB[18][26] ), .CI(\SUMB[18][27] ), 
        .CO(\CARRYB[19][26] ), .S(\SUMB[19][26] ) );
  FA_X1 S2_19_27 ( .A(\ab[19][27] ), .B(\CARRYB[18][27] ), .CI(\SUMB[18][28] ), 
        .CO(\CARRYB[19][27] ), .S(\SUMB[19][27] ) );
  FA_X1 S2_19_28 ( .A(\ab[19][28] ), .B(\CARRYB[18][28] ), .CI(\SUMB[18][29] ), 
        .CO(\CARRYB[19][28] ), .S(\SUMB[19][28] ) );
  FA_X1 S2_19_29 ( .A(\ab[19][29] ), .B(\CARRYB[18][29] ), .CI(\SUMB[18][30] ), 
        .CO(\CARRYB[19][29] ), .S(\SUMB[19][29] ) );
  FA_X1 S3_19_30 ( .A(\ab[19][30] ), .B(\CARRYB[18][30] ), .CI(\ab[18][31] ), 
        .CO(\CARRYB[19][30] ), .S(\SUMB[19][30] ) );
  FA_X1 S1_18_0 ( .A(\ab[18][0] ), .B(\CARRYB[17][0] ), .CI(\SUMB[17][1] ), 
        .CO(\CARRYB[18][0] ), .S(\A1[16] ) );
  FA_X1 S2_18_1 ( .A(\ab[18][1] ), .B(\CARRYB[17][1] ), .CI(\SUMB[17][2] ), 
        .CO(\CARRYB[18][1] ), .S(\SUMB[18][1] ) );
  FA_X1 S2_18_2 ( .A(\ab[18][2] ), .B(\CARRYB[17][2] ), .CI(\SUMB[17][3] ), 
        .CO(\CARRYB[18][2] ), .S(\SUMB[18][2] ) );
  FA_X1 S2_18_3 ( .A(\ab[18][3] ), .B(\CARRYB[17][3] ), .CI(\SUMB[17][4] ), 
        .CO(\CARRYB[18][3] ), .S(\SUMB[18][3] ) );
  FA_X1 S2_18_4 ( .A(\ab[18][4] ), .B(\CARRYB[17][4] ), .CI(\SUMB[17][5] ), 
        .CO(\CARRYB[18][4] ), .S(\SUMB[18][4] ) );
  FA_X1 S2_18_5 ( .A(\ab[18][5] ), .B(\CARRYB[17][5] ), .CI(\SUMB[17][6] ), 
        .CO(\CARRYB[18][5] ), .S(\SUMB[18][5] ) );
  FA_X1 S2_18_6 ( .A(\ab[18][6] ), .B(\CARRYB[17][6] ), .CI(\SUMB[17][7] ), 
        .CO(\CARRYB[18][6] ), .S(\SUMB[18][6] ) );
  FA_X1 S2_18_7 ( .A(\ab[18][7] ), .B(\CARRYB[17][7] ), .CI(\SUMB[17][8] ), 
        .CO(\CARRYB[18][7] ), .S(\SUMB[18][7] ) );
  FA_X1 S2_18_8 ( .A(\ab[18][8] ), .B(\CARRYB[17][8] ), .CI(\SUMB[17][9] ), 
        .CO(\CARRYB[18][8] ), .S(\SUMB[18][8] ) );
  FA_X1 S2_18_9 ( .A(\ab[18][9] ), .B(\CARRYB[17][9] ), .CI(\SUMB[17][10] ), 
        .CO(\CARRYB[18][9] ), .S(\SUMB[18][9] ) );
  FA_X1 S2_18_10 ( .A(\ab[18][10] ), .B(\CARRYB[17][10] ), .CI(\SUMB[17][11] ), 
        .CO(\CARRYB[18][10] ), .S(\SUMB[18][10] ) );
  FA_X1 S2_18_11 ( .A(\ab[18][11] ), .B(\CARRYB[17][11] ), .CI(\SUMB[17][12] ), 
        .CO(\CARRYB[18][11] ), .S(\SUMB[18][11] ) );
  FA_X1 S2_18_12 ( .A(\ab[18][12] ), .B(\CARRYB[17][12] ), .CI(\SUMB[17][13] ), 
        .CO(\CARRYB[18][12] ), .S(\SUMB[18][12] ) );
  FA_X1 S2_18_13 ( .A(\CARRYB[17][13] ), .B(\ab[18][13] ), .CI(\SUMB[17][14] ), 
        .CO(\CARRYB[18][13] ), .S(\SUMB[18][13] ) );
  FA_X1 S2_18_18 ( .A(\ab[18][18] ), .B(\CARRYB[17][18] ), .CI(\SUMB[17][19] ), 
        .CO(\CARRYB[18][18] ), .S(\SUMB[18][18] ) );
  FA_X1 S2_18_19 ( .A(\ab[18][19] ), .B(\CARRYB[17][19] ), .CI(\SUMB[17][20] ), 
        .CO(\CARRYB[18][19] ), .S(\SUMB[18][19] ) );
  FA_X1 S2_18_20 ( .A(\ab[18][20] ), .B(\CARRYB[17][20] ), .CI(\SUMB[17][21] ), 
        .CO(\CARRYB[18][20] ), .S(\SUMB[18][20] ) );
  FA_X1 S2_18_21 ( .A(\ab[18][21] ), .B(\CARRYB[17][21] ), .CI(\SUMB[17][22] ), 
        .CO(\CARRYB[18][21] ), .S(\SUMB[18][21] ) );
  FA_X1 S2_18_22 ( .A(\ab[18][22] ), .B(\CARRYB[17][22] ), .CI(\SUMB[17][23] ), 
        .CO(\CARRYB[18][22] ), .S(\SUMB[18][22] ) );
  FA_X1 S2_18_23 ( .A(\ab[18][23] ), .B(\CARRYB[17][23] ), .CI(\SUMB[17][24] ), 
        .CO(\CARRYB[18][23] ), .S(\SUMB[18][23] ) );
  FA_X1 S2_18_24 ( .A(\ab[18][24] ), .B(\CARRYB[17][24] ), .CI(\SUMB[17][25] ), 
        .CO(\CARRYB[18][24] ), .S(\SUMB[18][24] ) );
  FA_X1 S2_18_25 ( .A(\ab[18][25] ), .B(\CARRYB[17][25] ), .CI(\SUMB[17][26] ), 
        .CO(\CARRYB[18][25] ), .S(\SUMB[18][25] ) );
  FA_X1 S2_18_26 ( .A(\ab[18][26] ), .B(\CARRYB[17][26] ), .CI(\SUMB[17][27] ), 
        .CO(\CARRYB[18][26] ), .S(\SUMB[18][26] ) );
  FA_X1 S2_18_27 ( .A(\ab[18][27] ), .B(\CARRYB[17][27] ), .CI(\SUMB[17][28] ), 
        .CO(\CARRYB[18][27] ), .S(\SUMB[18][27] ) );
  FA_X1 S2_18_28 ( .A(\ab[18][28] ), .B(\CARRYB[17][28] ), .CI(\SUMB[17][29] ), 
        .CO(\CARRYB[18][28] ), .S(\SUMB[18][28] ) );
  FA_X1 S2_18_29 ( .A(\ab[18][29] ), .B(\CARRYB[17][29] ), .CI(\SUMB[17][30] ), 
        .CO(\CARRYB[18][29] ), .S(\SUMB[18][29] ) );
  FA_X1 S3_18_30 ( .A(\ab[18][30] ), .B(\CARRYB[17][30] ), .CI(\ab[17][31] ), 
        .CO(\CARRYB[18][30] ), .S(\SUMB[18][30] ) );
  FA_X1 S1_17_0 ( .A(\ab[17][0] ), .B(\CARRYB[16][0] ), .CI(\SUMB[16][1] ), 
        .CO(\CARRYB[17][0] ), .S(\A1[15] ) );
  FA_X1 S2_17_1 ( .A(\ab[17][1] ), .B(\CARRYB[16][1] ), .CI(\SUMB[16][2] ), 
        .CO(\CARRYB[17][1] ), .S(\SUMB[17][1] ) );
  FA_X1 S2_17_2 ( .A(\ab[17][2] ), .B(\CARRYB[16][2] ), .CI(\SUMB[16][3] ), 
        .CO(\CARRYB[17][2] ), .S(\SUMB[17][2] ) );
  FA_X1 S2_17_3 ( .A(\ab[17][3] ), .B(\CARRYB[16][3] ), .CI(\SUMB[16][4] ), 
        .CO(\CARRYB[17][3] ), .S(\SUMB[17][3] ) );
  FA_X1 S2_17_4 ( .A(\ab[17][4] ), .B(\CARRYB[16][4] ), .CI(\SUMB[16][5] ), 
        .CO(\CARRYB[17][4] ), .S(\SUMB[17][4] ) );
  FA_X1 S2_17_5 ( .A(\ab[17][5] ), .B(\CARRYB[16][5] ), .CI(\SUMB[16][6] ), 
        .CO(\CARRYB[17][5] ), .S(\SUMB[17][5] ) );
  FA_X1 S2_17_6 ( .A(\ab[17][6] ), .B(\CARRYB[16][6] ), .CI(\SUMB[16][7] ), 
        .CO(\CARRYB[17][6] ), .S(\SUMB[17][6] ) );
  FA_X1 S2_17_7 ( .A(\ab[17][7] ), .B(\CARRYB[16][7] ), .CI(\SUMB[16][8] ), 
        .CO(\CARRYB[17][7] ), .S(\SUMB[17][7] ) );
  FA_X1 S2_17_8 ( .A(\ab[17][8] ), .B(\CARRYB[16][8] ), .CI(\SUMB[16][9] ), 
        .CO(\CARRYB[17][8] ), .S(\SUMB[17][8] ) );
  FA_X1 S2_17_9 ( .A(\ab[17][9] ), .B(\CARRYB[16][9] ), .CI(\SUMB[16][10] ), 
        .CO(\CARRYB[17][9] ), .S(\SUMB[17][9] ) );
  FA_X1 S2_17_10 ( .A(\ab[17][10] ), .B(\CARRYB[16][10] ), .CI(\SUMB[16][11] ), 
        .CO(\CARRYB[17][10] ), .S(\SUMB[17][10] ) );
  FA_X1 S2_17_11 ( .A(\ab[17][11] ), .B(\CARRYB[16][11] ), .CI(\SUMB[16][12] ), 
        .CO(\CARRYB[17][11] ), .S(\SUMB[17][11] ) );
  FA_X1 S2_17_12 ( .A(\ab[17][12] ), .B(\CARRYB[16][12] ), .CI(\SUMB[16][13] ), 
        .CO(\CARRYB[17][12] ), .S(\SUMB[17][12] ) );
  FA_X1 S2_17_13 ( .A(\CARRYB[16][13] ), .B(\ab[17][13] ), .CI(\SUMB[16][14] ), 
        .CO(\CARRYB[17][13] ), .S(\SUMB[17][13] ) );
  FA_X1 S2_17_14 ( .A(\ab[17][14] ), .B(\CARRYB[16][14] ), .CI(\SUMB[16][15] ), 
        .CO(\CARRYB[17][14] ), .S(\SUMB[17][14] ) );
  FA_X1 S2_17_19 ( .A(\ab[17][19] ), .B(\CARRYB[16][19] ), .CI(\SUMB[16][20] ), 
        .CO(\CARRYB[17][19] ), .S(\SUMB[17][19] ) );
  FA_X1 S2_17_20 ( .A(\ab[17][20] ), .B(\CARRYB[16][20] ), .CI(\SUMB[16][21] ), 
        .CO(\CARRYB[17][20] ), .S(\SUMB[17][20] ) );
  FA_X1 S2_17_21 ( .A(\ab[17][21] ), .B(\CARRYB[16][21] ), .CI(\SUMB[16][22] ), 
        .CO(\CARRYB[17][21] ), .S(\SUMB[17][21] ) );
  FA_X1 S2_17_22 ( .A(\ab[17][22] ), .B(\CARRYB[16][22] ), .CI(\SUMB[16][23] ), 
        .CO(\CARRYB[17][22] ), .S(\SUMB[17][22] ) );
  FA_X1 S2_17_23 ( .A(\ab[17][23] ), .B(\CARRYB[16][23] ), .CI(\SUMB[16][24] ), 
        .CO(\CARRYB[17][23] ), .S(\SUMB[17][23] ) );
  FA_X1 S2_17_24 ( .A(\ab[17][24] ), .B(\CARRYB[16][24] ), .CI(\SUMB[16][25] ), 
        .CO(\CARRYB[17][24] ), .S(\SUMB[17][24] ) );
  FA_X1 S2_17_25 ( .A(\ab[17][25] ), .B(\CARRYB[16][25] ), .CI(\SUMB[16][26] ), 
        .CO(\CARRYB[17][25] ), .S(\SUMB[17][25] ) );
  FA_X1 S2_17_26 ( .A(\ab[17][26] ), .B(\CARRYB[16][26] ), .CI(\SUMB[16][27] ), 
        .CO(\CARRYB[17][26] ), .S(\SUMB[17][26] ) );
  FA_X1 S2_17_27 ( .A(\ab[17][27] ), .B(\CARRYB[16][27] ), .CI(\SUMB[16][28] ), 
        .CO(\CARRYB[17][27] ), .S(\SUMB[17][27] ) );
  FA_X1 S2_17_28 ( .A(\ab[17][28] ), .B(\CARRYB[16][28] ), .CI(\SUMB[16][29] ), 
        .CO(\CARRYB[17][28] ), .S(\SUMB[17][28] ) );
  FA_X1 S2_17_29 ( .A(\ab[17][29] ), .B(\CARRYB[16][29] ), .CI(\SUMB[16][30] ), 
        .CO(\CARRYB[17][29] ), .S(\SUMB[17][29] ) );
  FA_X1 S3_17_30 ( .A(\ab[17][30] ), .B(\CARRYB[16][30] ), .CI(\ab[16][31] ), 
        .CO(\CARRYB[17][30] ), .S(\SUMB[17][30] ) );
  FA_X1 S1_16_0 ( .A(\ab[16][0] ), .B(\CARRYB[15][0] ), .CI(\SUMB[15][1] ), 
        .CO(\CARRYB[16][0] ), .S(\A1[14] ) );
  FA_X1 S2_16_1 ( .A(\ab[16][1] ), .B(\CARRYB[15][1] ), .CI(\SUMB[15][2] ), 
        .CO(\CARRYB[16][1] ), .S(\SUMB[16][1] ) );
  FA_X1 S2_16_2 ( .A(\ab[16][2] ), .B(\CARRYB[15][2] ), .CI(\SUMB[15][3] ), 
        .CO(\CARRYB[16][2] ), .S(\SUMB[16][2] ) );
  FA_X1 S2_16_3 ( .A(\ab[16][3] ), .B(\CARRYB[15][3] ), .CI(\SUMB[15][4] ), 
        .CO(\CARRYB[16][3] ), .S(\SUMB[16][3] ) );
  FA_X1 S2_16_4 ( .A(\ab[16][4] ), .B(\CARRYB[15][4] ), .CI(\SUMB[15][5] ), 
        .CO(\CARRYB[16][4] ), .S(\SUMB[16][4] ) );
  FA_X1 S2_16_5 ( .A(\ab[16][5] ), .B(\CARRYB[15][5] ), .CI(\SUMB[15][6] ), 
        .CO(\CARRYB[16][5] ), .S(\SUMB[16][5] ) );
  FA_X1 S2_16_6 ( .A(\ab[16][6] ), .B(\CARRYB[15][6] ), .CI(\SUMB[15][7] ), 
        .CO(\CARRYB[16][6] ), .S(\SUMB[16][6] ) );
  FA_X1 S2_16_7 ( .A(\ab[16][7] ), .B(\CARRYB[15][7] ), .CI(\SUMB[15][8] ), 
        .CO(\CARRYB[16][7] ), .S(\SUMB[16][7] ) );
  FA_X1 S2_16_8 ( .A(\ab[16][8] ), .B(\CARRYB[15][8] ), .CI(\SUMB[15][9] ), 
        .CO(\CARRYB[16][8] ), .S(\SUMB[16][8] ) );
  FA_X1 S2_16_9 ( .A(\ab[16][9] ), .B(\CARRYB[15][9] ), .CI(\SUMB[15][10] ), 
        .CO(\CARRYB[16][9] ), .S(\SUMB[16][9] ) );
  FA_X1 S2_16_10 ( .A(\ab[16][10] ), .B(\CARRYB[15][10] ), .CI(\SUMB[15][11] ), 
        .CO(\CARRYB[16][10] ), .S(\SUMB[16][10] ) );
  FA_X1 S2_16_11 ( .A(\ab[16][11] ), .B(\CARRYB[15][11] ), .CI(\SUMB[15][12] ), 
        .CO(\CARRYB[16][11] ), .S(\SUMB[16][11] ) );
  FA_X1 S2_16_12 ( .A(\ab[16][12] ), .B(\CARRYB[15][12] ), .CI(\SUMB[15][13] ), 
        .CO(\CARRYB[16][12] ), .S(\SUMB[16][12] ) );
  FA_X1 S2_16_13 ( .A(\ab[16][13] ), .B(\CARRYB[15][13] ), .CI(\SUMB[15][14] ), 
        .CO(\CARRYB[16][13] ), .S(\SUMB[16][13] ) );
  FA_X1 S2_16_14 ( .A(\ab[16][14] ), .B(\CARRYB[15][14] ), .CI(\SUMB[15][15] ), 
        .CO(\CARRYB[16][14] ), .S(\SUMB[16][14] ) );
  FA_X1 S2_16_15 ( .A(\ab[16][15] ), .B(\CARRYB[15][15] ), .CI(\SUMB[15][16] ), 
        .CO(\CARRYB[16][15] ), .S(\SUMB[16][15] ) );
  FA_X1 S2_16_20 ( .A(\ab[16][20] ), .B(\CARRYB[15][20] ), .CI(\SUMB[15][21] ), 
        .CO(\CARRYB[16][20] ), .S(\SUMB[16][20] ) );
  FA_X1 S2_16_21 ( .A(\ab[16][21] ), .B(\CARRYB[15][21] ), .CI(\SUMB[15][22] ), 
        .CO(\CARRYB[16][21] ), .S(\SUMB[16][21] ) );
  FA_X1 S2_16_22 ( .A(\ab[16][22] ), .B(\CARRYB[15][22] ), .CI(\SUMB[15][23] ), 
        .CO(\CARRYB[16][22] ), .S(\SUMB[16][22] ) );
  FA_X1 S2_16_23 ( .A(\ab[16][23] ), .B(\CARRYB[15][23] ), .CI(\SUMB[15][24] ), 
        .CO(\CARRYB[16][23] ), .S(\SUMB[16][23] ) );
  FA_X1 S2_16_24 ( .A(\ab[16][24] ), .B(\CARRYB[15][24] ), .CI(\SUMB[15][25] ), 
        .CO(\CARRYB[16][24] ), .S(\SUMB[16][24] ) );
  FA_X1 S2_16_25 ( .A(\ab[16][25] ), .B(\CARRYB[15][25] ), .CI(\SUMB[15][26] ), 
        .CO(\CARRYB[16][25] ), .S(\SUMB[16][25] ) );
  FA_X1 S2_16_26 ( .A(\ab[16][26] ), .B(\CARRYB[15][26] ), .CI(\SUMB[15][27] ), 
        .CO(\CARRYB[16][26] ), .S(\SUMB[16][26] ) );
  FA_X1 S2_16_27 ( .A(\ab[16][27] ), .B(\CARRYB[15][27] ), .CI(\SUMB[15][28] ), 
        .CO(\CARRYB[16][27] ), .S(\SUMB[16][27] ) );
  FA_X1 S2_16_28 ( .A(\ab[16][28] ), .B(\CARRYB[15][28] ), .CI(\SUMB[15][29] ), 
        .CO(\CARRYB[16][28] ), .S(\SUMB[16][28] ) );
  FA_X1 S2_16_29 ( .A(\ab[16][29] ), .B(\CARRYB[15][29] ), .CI(\SUMB[15][30] ), 
        .CO(\CARRYB[16][29] ), .S(\SUMB[16][29] ) );
  FA_X1 S3_16_30 ( .A(\ab[16][30] ), .B(\CARRYB[15][30] ), .CI(\ab[15][31] ), 
        .CO(\CARRYB[16][30] ), .S(\SUMB[16][30] ) );
  FA_X1 S1_15_0 ( .A(\ab[15][0] ), .B(\CARRYB[14][0] ), .CI(\SUMB[14][1] ), 
        .CO(\CARRYB[15][0] ), .S(\A1[13] ) );
  FA_X1 S2_15_1 ( .A(\ab[15][1] ), .B(\CARRYB[14][1] ), .CI(\SUMB[14][2] ), 
        .CO(\CARRYB[15][1] ), .S(\SUMB[15][1] ) );
  FA_X1 S2_15_2 ( .A(\ab[15][2] ), .B(\CARRYB[14][2] ), .CI(\SUMB[14][3] ), 
        .CO(\CARRYB[15][2] ), .S(\SUMB[15][2] ) );
  FA_X1 S2_15_3 ( .A(\ab[15][3] ), .B(\CARRYB[14][3] ), .CI(\SUMB[14][4] ), 
        .CO(\CARRYB[15][3] ), .S(\SUMB[15][3] ) );
  FA_X1 S2_15_4 ( .A(\ab[15][4] ), .B(\CARRYB[14][4] ), .CI(\SUMB[14][5] ), 
        .CO(\CARRYB[15][4] ), .S(\SUMB[15][4] ) );
  FA_X1 S2_15_5 ( .A(\ab[15][5] ), .B(\CARRYB[14][5] ), .CI(\SUMB[14][6] ), 
        .CO(\CARRYB[15][5] ), .S(\SUMB[15][5] ) );
  FA_X1 S2_15_6 ( .A(\ab[15][6] ), .B(\CARRYB[14][6] ), .CI(\SUMB[14][7] ), 
        .CO(\CARRYB[15][6] ), .S(\SUMB[15][6] ) );
  FA_X1 S2_15_7 ( .A(\ab[15][7] ), .B(\CARRYB[14][7] ), .CI(\SUMB[14][8] ), 
        .CO(\CARRYB[15][7] ), .S(\SUMB[15][7] ) );
  FA_X1 S2_15_8 ( .A(\ab[15][8] ), .B(\CARRYB[14][8] ), .CI(\SUMB[14][9] ), 
        .CO(\CARRYB[15][8] ), .S(\SUMB[15][8] ) );
  FA_X1 S2_15_9 ( .A(\ab[15][9] ), .B(\CARRYB[14][9] ), .CI(\SUMB[14][10] ), 
        .CO(\CARRYB[15][9] ), .S(\SUMB[15][9] ) );
  FA_X1 S2_15_10 ( .A(\ab[15][10] ), .B(\CARRYB[14][10] ), .CI(\SUMB[14][11] ), 
        .CO(\CARRYB[15][10] ), .S(\SUMB[15][10] ) );
  FA_X1 S2_15_11 ( .A(\ab[15][11] ), .B(\CARRYB[14][11] ), .CI(\SUMB[14][12] ), 
        .CO(\CARRYB[15][11] ), .S(\SUMB[15][11] ) );
  FA_X1 S2_15_12 ( .A(\ab[15][12] ), .B(\CARRYB[14][12] ), .CI(\SUMB[14][13] ), 
        .CO(\CARRYB[15][12] ), .S(\SUMB[15][12] ) );
  FA_X1 S2_15_13 ( .A(\ab[15][13] ), .B(\CARRYB[14][13] ), .CI(\SUMB[14][14] ), 
        .CO(\CARRYB[15][13] ), .S(\SUMB[15][13] ) );
  FA_X1 S2_15_14 ( .A(\ab[15][14] ), .B(\CARRYB[14][14] ), .CI(\SUMB[14][15] ), 
        .CO(\CARRYB[15][14] ), .S(\SUMB[15][14] ) );
  FA_X1 S2_15_15 ( .A(\ab[15][15] ), .B(\CARRYB[14][15] ), .CI(\SUMB[14][16] ), 
        .CO(\CARRYB[15][15] ), .S(\SUMB[15][15] ) );
  FA_X1 S2_15_16 ( .A(\ab[15][16] ), .B(\CARRYB[14][16] ), .CI(\SUMB[14][17] ), 
        .CO(\CARRYB[15][16] ), .S(\SUMB[15][16] ) );
  FA_X1 S2_15_21 ( .A(\ab[15][21] ), .B(\CARRYB[14][21] ), .CI(\SUMB[14][22] ), 
        .CO(\CARRYB[15][21] ), .S(\SUMB[15][21] ) );
  FA_X1 S2_15_22 ( .A(\ab[15][22] ), .B(\CARRYB[14][22] ), .CI(\SUMB[14][23] ), 
        .CO(\CARRYB[15][22] ), .S(\SUMB[15][22] ) );
  FA_X1 S2_15_23 ( .A(\ab[15][23] ), .B(\CARRYB[14][23] ), .CI(\SUMB[14][24] ), 
        .CO(\CARRYB[15][23] ), .S(\SUMB[15][23] ) );
  FA_X1 S2_15_24 ( .A(\ab[15][24] ), .B(\CARRYB[14][24] ), .CI(\SUMB[14][25] ), 
        .CO(\CARRYB[15][24] ), .S(\SUMB[15][24] ) );
  FA_X1 S2_15_25 ( .A(\ab[15][25] ), .B(\CARRYB[14][25] ), .CI(\SUMB[14][26] ), 
        .CO(\CARRYB[15][25] ), .S(\SUMB[15][25] ) );
  FA_X1 S2_15_26 ( .A(\ab[15][26] ), .B(\CARRYB[14][26] ), .CI(\SUMB[14][27] ), 
        .CO(\CARRYB[15][26] ), .S(\SUMB[15][26] ) );
  FA_X1 S2_15_27 ( .A(\ab[15][27] ), .B(\CARRYB[14][27] ), .CI(\SUMB[14][28] ), 
        .CO(\CARRYB[15][27] ), .S(\SUMB[15][27] ) );
  FA_X1 S2_15_28 ( .A(\ab[15][28] ), .B(\CARRYB[14][28] ), .CI(\SUMB[14][29] ), 
        .CO(\CARRYB[15][28] ), .S(\SUMB[15][28] ) );
  FA_X1 S2_15_29 ( .A(\ab[15][29] ), .B(\CARRYB[14][29] ), .CI(\SUMB[14][30] ), 
        .CO(\CARRYB[15][29] ), .S(\SUMB[15][29] ) );
  FA_X1 S3_15_30 ( .A(\ab[15][30] ), .B(\CARRYB[14][30] ), .CI(\ab[14][31] ), 
        .CO(\CARRYB[15][30] ), .S(\SUMB[15][30] ) );
  FA_X1 S1_14_0 ( .A(\ab[14][0] ), .B(\CARRYB[13][0] ), .CI(\SUMB[13][1] ), 
        .CO(\CARRYB[14][0] ), .S(\A1[12] ) );
  FA_X1 S2_14_1 ( .A(\ab[14][1] ), .B(\CARRYB[13][1] ), .CI(\SUMB[13][2] ), 
        .CO(\CARRYB[14][1] ), .S(\SUMB[14][1] ) );
  FA_X1 S2_14_2 ( .A(\ab[14][2] ), .B(\CARRYB[13][2] ), .CI(\SUMB[13][3] ), 
        .CO(\CARRYB[14][2] ), .S(\SUMB[14][2] ) );
  FA_X1 S2_14_3 ( .A(\ab[14][3] ), .B(\CARRYB[13][3] ), .CI(\SUMB[13][4] ), 
        .CO(\CARRYB[14][3] ), .S(\SUMB[14][3] ) );
  FA_X1 S2_14_4 ( .A(\ab[14][4] ), .B(\CARRYB[13][4] ), .CI(\SUMB[13][5] ), 
        .CO(\CARRYB[14][4] ), .S(\SUMB[14][4] ) );
  FA_X1 S2_14_5 ( .A(\ab[14][5] ), .B(\CARRYB[13][5] ), .CI(\SUMB[13][6] ), 
        .CO(\CARRYB[14][5] ), .S(\SUMB[14][5] ) );
  FA_X1 S2_14_6 ( .A(\ab[14][6] ), .B(\CARRYB[13][6] ), .CI(\SUMB[13][7] ), 
        .CO(\CARRYB[14][6] ), .S(\SUMB[14][6] ) );
  FA_X1 S2_14_7 ( .A(\ab[14][7] ), .B(\CARRYB[13][7] ), .CI(\SUMB[13][8] ), 
        .CO(\CARRYB[14][7] ), .S(\SUMB[14][7] ) );
  FA_X1 S2_14_8 ( .A(\ab[14][8] ), .B(\CARRYB[13][8] ), .CI(\SUMB[13][9] ), 
        .CO(\CARRYB[14][8] ), .S(\SUMB[14][8] ) );
  FA_X1 S2_14_9 ( .A(\ab[14][9] ), .B(\CARRYB[13][9] ), .CI(\SUMB[13][10] ), 
        .CO(\CARRYB[14][9] ), .S(\SUMB[14][9] ) );
  FA_X1 S2_14_10 ( .A(\ab[14][10] ), .B(\CARRYB[13][10] ), .CI(\SUMB[13][11] ), 
        .CO(\CARRYB[14][10] ), .S(\SUMB[14][10] ) );
  FA_X1 S2_14_11 ( .A(\ab[14][11] ), .B(\CARRYB[13][11] ), .CI(\SUMB[13][12] ), 
        .CO(\CARRYB[14][11] ), .S(\SUMB[14][11] ) );
  FA_X1 S2_14_12 ( .A(\ab[14][12] ), .B(\CARRYB[13][12] ), .CI(\SUMB[13][13] ), 
        .CO(\CARRYB[14][12] ), .S(\SUMB[14][12] ) );
  FA_X1 S2_14_13 ( .A(\ab[14][13] ), .B(\CARRYB[13][13] ), .CI(\SUMB[13][14] ), 
        .CO(\CARRYB[14][13] ), .S(\SUMB[14][13] ) );
  FA_X1 S2_14_14 ( .A(\ab[14][14] ), .B(\CARRYB[13][14] ), .CI(\SUMB[13][15] ), 
        .CO(\CARRYB[14][14] ), .S(\SUMB[14][14] ) );
  FA_X1 S2_14_15 ( .A(\ab[14][15] ), .B(\CARRYB[13][15] ), .CI(\SUMB[13][16] ), 
        .CO(\CARRYB[14][15] ), .S(\SUMB[14][15] ) );
  FA_X1 S2_14_16 ( .A(\ab[14][16] ), .B(\CARRYB[13][16] ), .CI(\SUMB[13][17] ), 
        .CO(\CARRYB[14][16] ), .S(\SUMB[14][16] ) );
  FA_X1 S2_14_17 ( .A(\CARRYB[13][17] ), .B(\ab[14][17] ), .CI(\SUMB[13][18] ), 
        .CO(\CARRYB[14][17] ), .S(\SUMB[14][17] ) );
  FA_X1 S2_14_22 ( .A(\ab[14][22] ), .B(\CARRYB[13][22] ), .CI(\SUMB[13][23] ), 
        .CO(\CARRYB[14][22] ), .S(\SUMB[14][22] ) );
  FA_X1 S2_14_23 ( .A(\ab[14][23] ), .B(\CARRYB[13][23] ), .CI(\SUMB[13][24] ), 
        .CO(\CARRYB[14][23] ), .S(\SUMB[14][23] ) );
  FA_X1 S2_14_24 ( .A(\ab[14][24] ), .B(\CARRYB[13][24] ), .CI(\SUMB[13][25] ), 
        .CO(\CARRYB[14][24] ), .S(\SUMB[14][24] ) );
  FA_X1 S2_14_25 ( .A(\ab[14][25] ), .B(\CARRYB[13][25] ), .CI(\SUMB[13][26] ), 
        .CO(\CARRYB[14][25] ), .S(\SUMB[14][25] ) );
  FA_X1 S2_14_26 ( .A(\ab[14][26] ), .B(\CARRYB[13][26] ), .CI(\SUMB[13][27] ), 
        .CO(\CARRYB[14][26] ), .S(\SUMB[14][26] ) );
  FA_X1 S2_14_27 ( .A(\ab[14][27] ), .B(\CARRYB[13][27] ), .CI(\SUMB[13][28] ), 
        .CO(\CARRYB[14][27] ), .S(\SUMB[14][27] ) );
  FA_X1 S2_14_28 ( .A(\ab[14][28] ), .B(\CARRYB[13][28] ), .CI(\SUMB[13][29] ), 
        .CO(\CARRYB[14][28] ), .S(\SUMB[14][28] ) );
  FA_X1 S2_14_29 ( .A(\ab[14][29] ), .B(\CARRYB[13][29] ), .CI(\SUMB[13][30] ), 
        .CO(\CARRYB[14][29] ), .S(\SUMB[14][29] ) );
  FA_X1 S3_14_30 ( .A(\ab[14][30] ), .B(\CARRYB[13][30] ), .CI(\ab[13][31] ), 
        .CO(\CARRYB[14][30] ), .S(\SUMB[14][30] ) );
  FA_X1 S1_13_0 ( .A(\ab[13][0] ), .B(\CARRYB[12][0] ), .CI(\SUMB[12][1] ), 
        .CO(\CARRYB[13][0] ), .S(\A1[11] ) );
  FA_X1 S2_13_1 ( .A(\ab[13][1] ), .B(\CARRYB[12][1] ), .CI(\SUMB[12][2] ), 
        .CO(\CARRYB[13][1] ), .S(\SUMB[13][1] ) );
  FA_X1 S2_13_2 ( .A(\ab[13][2] ), .B(\CARRYB[12][2] ), .CI(\SUMB[12][3] ), 
        .CO(\CARRYB[13][2] ), .S(\SUMB[13][2] ) );
  FA_X1 S2_13_3 ( .A(\ab[13][3] ), .B(\CARRYB[12][3] ), .CI(\SUMB[12][4] ), 
        .CO(\CARRYB[13][3] ), .S(\SUMB[13][3] ) );
  FA_X1 S2_13_4 ( .A(\ab[13][4] ), .B(\CARRYB[12][4] ), .CI(\SUMB[12][5] ), 
        .CO(\CARRYB[13][4] ), .S(\SUMB[13][4] ) );
  FA_X1 S2_13_5 ( .A(\ab[13][5] ), .B(\CARRYB[12][5] ), .CI(\SUMB[12][6] ), 
        .CO(\CARRYB[13][5] ), .S(\SUMB[13][5] ) );
  FA_X1 S2_13_6 ( .A(\ab[13][6] ), .B(\CARRYB[12][6] ), .CI(\SUMB[12][7] ), 
        .CO(\CARRYB[13][6] ), .S(\SUMB[13][6] ) );
  FA_X1 S2_13_7 ( .A(\ab[13][7] ), .B(\CARRYB[12][7] ), .CI(\SUMB[12][8] ), 
        .CO(\CARRYB[13][7] ), .S(\SUMB[13][7] ) );
  FA_X1 S2_13_8 ( .A(\ab[13][8] ), .B(\CARRYB[12][8] ), .CI(\SUMB[12][9] ), 
        .CO(\CARRYB[13][8] ), .S(\SUMB[13][8] ) );
  FA_X1 S2_13_9 ( .A(\ab[13][9] ), .B(\CARRYB[12][9] ), .CI(\SUMB[12][10] ), 
        .CO(\CARRYB[13][9] ), .S(\SUMB[13][9] ) );
  FA_X1 S2_13_10 ( .A(\ab[13][10] ), .B(\CARRYB[12][10] ), .CI(\SUMB[12][11] ), 
        .CO(\CARRYB[13][10] ), .S(\SUMB[13][10] ) );
  FA_X1 S2_13_11 ( .A(\ab[13][11] ), .B(\CARRYB[12][11] ), .CI(\SUMB[12][12] ), 
        .CO(\CARRYB[13][11] ), .S(\SUMB[13][11] ) );
  FA_X1 S2_13_12 ( .A(\ab[13][12] ), .B(\CARRYB[12][12] ), .CI(\SUMB[12][13] ), 
        .CO(\CARRYB[13][12] ), .S(\SUMB[13][12] ) );
  FA_X1 S2_13_13 ( .A(\ab[13][13] ), .B(\CARRYB[12][13] ), .CI(\SUMB[12][14] ), 
        .CO(\CARRYB[13][13] ), .S(\SUMB[13][13] ) );
  FA_X1 S2_13_14 ( .A(\ab[13][14] ), .B(\CARRYB[12][14] ), .CI(\SUMB[12][15] ), 
        .CO(\CARRYB[13][14] ), .S(\SUMB[13][14] ) );
  FA_X1 S2_13_15 ( .A(\CARRYB[12][15] ), .B(\ab[13][15] ), .CI(\SUMB[12][16] ), 
        .CO(\CARRYB[13][15] ), .S(\SUMB[13][15] ) );
  FA_X1 S2_13_16 ( .A(\ab[13][16] ), .B(\CARRYB[12][16] ), .CI(\SUMB[12][17] ), 
        .CO(\CARRYB[13][16] ), .S(\SUMB[13][16] ) );
  FA_X1 S2_13_17 ( .A(\CARRYB[12][17] ), .B(\ab[13][17] ), .CI(\SUMB[12][18] ), 
        .CO(\CARRYB[13][17] ), .S(\SUMB[13][17] ) );
  FA_X1 S2_13_18 ( .A(\ab[13][18] ), .B(\CARRYB[12][18] ), .CI(\SUMB[12][19] ), 
        .CO(\CARRYB[13][18] ), .S(\SUMB[13][18] ) );
  FA_X1 S2_13_23 ( .A(\ab[13][23] ), .B(\CARRYB[12][23] ), .CI(\SUMB[12][24] ), 
        .CO(\CARRYB[13][23] ), .S(\SUMB[13][23] ) );
  FA_X1 S2_13_24 ( .A(\ab[13][24] ), .B(\CARRYB[12][24] ), .CI(\SUMB[12][25] ), 
        .CO(\CARRYB[13][24] ), .S(\SUMB[13][24] ) );
  FA_X1 S2_13_25 ( .A(\ab[13][25] ), .B(\CARRYB[12][25] ), .CI(\SUMB[12][26] ), 
        .CO(\CARRYB[13][25] ), .S(\SUMB[13][25] ) );
  FA_X1 S2_13_26 ( .A(\ab[13][26] ), .B(\CARRYB[12][26] ), .CI(\SUMB[12][27] ), 
        .CO(\CARRYB[13][26] ), .S(\SUMB[13][26] ) );
  FA_X1 S2_13_27 ( .A(\ab[13][27] ), .B(\CARRYB[12][27] ), .CI(\SUMB[12][28] ), 
        .CO(\CARRYB[13][27] ), .S(\SUMB[13][27] ) );
  FA_X1 S2_13_28 ( .A(\ab[13][28] ), .B(\CARRYB[12][28] ), .CI(\SUMB[12][29] ), 
        .CO(\CARRYB[13][28] ), .S(\SUMB[13][28] ) );
  FA_X1 S2_13_29 ( .A(\ab[13][29] ), .B(\CARRYB[12][29] ), .CI(\SUMB[12][30] ), 
        .CO(\CARRYB[13][29] ), .S(\SUMB[13][29] ) );
  FA_X1 S3_13_30 ( .A(\ab[13][30] ), .B(\CARRYB[12][30] ), .CI(\ab[12][31] ), 
        .CO(\CARRYB[13][30] ), .S(\SUMB[13][30] ) );
  FA_X1 S1_12_0 ( .A(\ab[12][0] ), .B(\CARRYB[11][0] ), .CI(\SUMB[11][1] ), 
        .CO(\CARRYB[12][0] ), .S(\A1[10] ) );
  FA_X1 S2_12_1 ( .A(\ab[12][1] ), .B(\CARRYB[11][1] ), .CI(\SUMB[11][2] ), 
        .CO(\CARRYB[12][1] ), .S(\SUMB[12][1] ) );
  FA_X1 S2_12_2 ( .A(\ab[12][2] ), .B(\CARRYB[11][2] ), .CI(\SUMB[11][3] ), 
        .CO(\CARRYB[12][2] ), .S(\SUMB[12][2] ) );
  FA_X1 S2_12_3 ( .A(\ab[12][3] ), .B(\CARRYB[11][3] ), .CI(\SUMB[11][4] ), 
        .CO(\CARRYB[12][3] ), .S(\SUMB[12][3] ) );
  FA_X1 S2_12_4 ( .A(\ab[12][4] ), .B(\CARRYB[11][4] ), .CI(\SUMB[11][5] ), 
        .CO(\CARRYB[12][4] ), .S(\SUMB[12][4] ) );
  FA_X1 S2_12_5 ( .A(\ab[12][5] ), .B(\CARRYB[11][5] ), .CI(\SUMB[11][6] ), 
        .CO(\CARRYB[12][5] ), .S(\SUMB[12][5] ) );
  FA_X1 S2_12_6 ( .A(\ab[12][6] ), .B(\CARRYB[11][6] ), .CI(\SUMB[11][7] ), 
        .CO(\CARRYB[12][6] ), .S(\SUMB[12][6] ) );
  FA_X1 S2_12_7 ( .A(\ab[12][7] ), .B(\CARRYB[11][7] ), .CI(\SUMB[11][8] ), 
        .CO(\CARRYB[12][7] ), .S(\SUMB[12][7] ) );
  FA_X1 S2_12_8 ( .A(\ab[12][8] ), .B(\CARRYB[11][8] ), .CI(\SUMB[11][9] ), 
        .CO(\CARRYB[12][8] ), .S(\SUMB[12][8] ) );
  FA_X1 S2_12_9 ( .A(\ab[12][9] ), .B(\CARRYB[11][9] ), .CI(\SUMB[11][10] ), 
        .CO(\CARRYB[12][9] ), .S(\SUMB[12][9] ) );
  FA_X1 S2_12_10 ( .A(\ab[12][10] ), .B(\CARRYB[11][10] ), .CI(\SUMB[11][11] ), 
        .CO(\CARRYB[12][10] ), .S(\SUMB[12][10] ) );
  FA_X1 S2_12_11 ( .A(\ab[12][11] ), .B(\CARRYB[11][11] ), .CI(\SUMB[11][12] ), 
        .CO(\CARRYB[12][11] ), .S(\SUMB[12][11] ) );
  FA_X1 S2_12_12 ( .A(\ab[12][12] ), .B(\CARRYB[11][12] ), .CI(\SUMB[11][13] ), 
        .CO(\CARRYB[12][12] ), .S(\SUMB[12][12] ) );
  FA_X1 S2_12_13 ( .A(\ab[12][13] ), .B(\CARRYB[11][13] ), .CI(\SUMB[11][14] ), 
        .CO(\CARRYB[12][13] ), .S(\SUMB[12][13] ) );
  FA_X1 S2_12_14 ( .A(\ab[12][14] ), .B(\CARRYB[11][14] ), .CI(\SUMB[11][15] ), 
        .CO(\CARRYB[12][14] ), .S(\SUMB[12][14] ) );
  FA_X1 S2_12_15 ( .A(\ab[12][15] ), .B(\CARRYB[11][15] ), .CI(\SUMB[11][16] ), 
        .CO(\CARRYB[12][15] ), .S(\SUMB[12][15] ) );
  FA_X1 S2_12_16 ( .A(\ab[12][16] ), .B(\CARRYB[11][16] ), .CI(\SUMB[11][17] ), 
        .CO(\CARRYB[12][16] ), .S(\SUMB[12][16] ) );
  FA_X1 S2_12_17 ( .A(\ab[12][17] ), .B(\CARRYB[11][17] ), .CI(\SUMB[11][18] ), 
        .CO(\CARRYB[12][17] ), .S(\SUMB[12][17] ) );
  FA_X1 S2_12_18 ( .A(\CARRYB[11][18] ), .B(\ab[12][18] ), .CI(\SUMB[11][19] ), 
        .CO(\CARRYB[12][18] ), .S(\SUMB[12][18] ) );
  FA_X1 S2_12_19 ( .A(\CARRYB[11][19] ), .B(\ab[12][19] ), .CI(\SUMB[11][20] ), 
        .CO(\CARRYB[12][19] ), .S(\SUMB[12][19] ) );
  FA_X1 S2_12_24 ( .A(\ab[12][24] ), .B(\CARRYB[11][24] ), .CI(\SUMB[11][25] ), 
        .CO(\CARRYB[12][24] ), .S(\SUMB[12][24] ) );
  FA_X1 S2_12_25 ( .A(\ab[12][25] ), .B(\CARRYB[11][25] ), .CI(\SUMB[11][26] ), 
        .CO(\CARRYB[12][25] ), .S(\SUMB[12][25] ) );
  FA_X1 S2_12_26 ( .A(\ab[12][26] ), .B(\CARRYB[11][26] ), .CI(\SUMB[11][27] ), 
        .CO(\CARRYB[12][26] ), .S(\SUMB[12][26] ) );
  FA_X1 S2_12_27 ( .A(\ab[12][27] ), .B(\CARRYB[11][27] ), .CI(\SUMB[11][28] ), 
        .CO(\CARRYB[12][27] ), .S(\SUMB[12][27] ) );
  FA_X1 S2_12_28 ( .A(\ab[12][28] ), .B(\CARRYB[11][28] ), .CI(\SUMB[11][29] ), 
        .CO(\CARRYB[12][28] ), .S(\SUMB[12][28] ) );
  FA_X1 S2_12_29 ( .A(\ab[12][29] ), .B(\CARRYB[11][29] ), .CI(\SUMB[11][30] ), 
        .CO(\CARRYB[12][29] ), .S(\SUMB[12][29] ) );
  FA_X1 S3_12_30 ( .A(\ab[12][30] ), .B(\CARRYB[11][30] ), .CI(\ab[11][31] ), 
        .CO(\CARRYB[12][30] ), .S(\SUMB[12][30] ) );
  FA_X1 S1_11_0 ( .A(\ab[11][0] ), .B(\CARRYB[10][0] ), .CI(\SUMB[10][1] ), 
        .CO(\CARRYB[11][0] ), .S(\A1[9] ) );
  FA_X1 S2_11_1 ( .A(\ab[11][1] ), .B(\CARRYB[10][1] ), .CI(\SUMB[10][2] ), 
        .CO(\CARRYB[11][1] ), .S(\SUMB[11][1] ) );
  FA_X1 S2_11_2 ( .A(\ab[11][2] ), .B(\CARRYB[10][2] ), .CI(\SUMB[10][3] ), 
        .CO(\CARRYB[11][2] ), .S(\SUMB[11][2] ) );
  FA_X1 S2_11_3 ( .A(\ab[11][3] ), .B(\CARRYB[10][3] ), .CI(\SUMB[10][4] ), 
        .CO(\CARRYB[11][3] ), .S(\SUMB[11][3] ) );
  FA_X1 S2_11_4 ( .A(\ab[11][4] ), .B(\CARRYB[10][4] ), .CI(\SUMB[10][5] ), 
        .CO(\CARRYB[11][4] ), .S(\SUMB[11][4] ) );
  FA_X1 S2_11_5 ( .A(\ab[11][5] ), .B(\CARRYB[10][5] ), .CI(\SUMB[10][6] ), 
        .CO(\CARRYB[11][5] ), .S(\SUMB[11][5] ) );
  FA_X1 S2_11_6 ( .A(\ab[11][6] ), .B(\CARRYB[10][6] ), .CI(\SUMB[10][7] ), 
        .CO(\CARRYB[11][6] ), .S(\SUMB[11][6] ) );
  FA_X1 S2_11_7 ( .A(\ab[11][7] ), .B(\CARRYB[10][7] ), .CI(\SUMB[10][8] ), 
        .CO(\CARRYB[11][7] ), .S(\SUMB[11][7] ) );
  FA_X1 S2_11_8 ( .A(\ab[11][8] ), .B(\CARRYB[10][8] ), .CI(\SUMB[10][9] ), 
        .CO(\CARRYB[11][8] ), .S(\SUMB[11][8] ) );
  FA_X1 S2_11_9 ( .A(\ab[11][9] ), .B(\CARRYB[10][9] ), .CI(\SUMB[10][10] ), 
        .CO(\CARRYB[11][9] ), .S(\SUMB[11][9] ) );
  FA_X1 S2_11_10 ( .A(\ab[11][10] ), .B(\CARRYB[10][10] ), .CI(\SUMB[10][11] ), 
        .CO(\CARRYB[11][10] ), .S(\SUMB[11][10] ) );
  FA_X1 S2_11_11 ( .A(\ab[11][11] ), .B(\CARRYB[10][11] ), .CI(\SUMB[10][12] ), 
        .CO(\CARRYB[11][11] ), .S(\SUMB[11][11] ) );
  FA_X1 S2_11_12 ( .A(\ab[11][12] ), .B(\CARRYB[10][12] ), .CI(\SUMB[10][13] ), 
        .CO(\CARRYB[11][12] ), .S(\SUMB[11][12] ) );
  FA_X1 S2_11_13 ( .A(\ab[11][13] ), .B(\CARRYB[10][13] ), .CI(\SUMB[10][14] ), 
        .CO(\CARRYB[11][13] ), .S(\SUMB[11][13] ) );
  FA_X1 S2_11_14 ( .A(\ab[11][14] ), .B(\CARRYB[10][14] ), .CI(\SUMB[10][15] ), 
        .CO(\CARRYB[11][14] ), .S(\SUMB[11][14] ) );
  FA_X1 S2_11_15 ( .A(\ab[11][15] ), .B(\CARRYB[10][15] ), .CI(\SUMB[10][16] ), 
        .CO(\CARRYB[11][15] ), .S(\SUMB[11][15] ) );
  FA_X1 S2_11_16 ( .A(\ab[11][16] ), .B(\CARRYB[10][16] ), .CI(\SUMB[10][17] ), 
        .CO(\CARRYB[11][16] ), .S(\SUMB[11][16] ) );
  FA_X1 S2_11_17 ( .A(\ab[11][17] ), .B(\CARRYB[10][17] ), .CI(\SUMB[10][18] ), 
        .CO(\CARRYB[11][17] ), .S(\SUMB[11][17] ) );
  FA_X1 S2_11_18 ( .A(\ab[11][18] ), .B(\CARRYB[10][18] ), .CI(\SUMB[10][19] ), 
        .CO(\CARRYB[11][18] ), .S(\SUMB[11][18] ) );
  FA_X1 S2_11_19 ( .A(\CARRYB[10][19] ), .B(\ab[11][19] ), .CI(\SUMB[10][20] ), 
        .CO(\CARRYB[11][19] ), .S(\SUMB[11][19] ) );
  FA_X1 S2_11_20 ( .A(\ab[11][20] ), .B(\CARRYB[10][20] ), .CI(\SUMB[10][21] ), 
        .CO(\CARRYB[11][20] ), .S(\SUMB[11][20] ) );
  FA_X1 S2_11_25 ( .A(\ab[11][25] ), .B(\CARRYB[10][25] ), .CI(\SUMB[10][26] ), 
        .CO(\CARRYB[11][25] ), .S(\SUMB[11][25] ) );
  FA_X1 S2_11_26 ( .A(\ab[11][26] ), .B(\CARRYB[10][26] ), .CI(\SUMB[10][27] ), 
        .CO(\CARRYB[11][26] ), .S(\SUMB[11][26] ) );
  FA_X1 S2_11_27 ( .A(\ab[11][27] ), .B(\CARRYB[10][27] ), .CI(\SUMB[10][28] ), 
        .CO(\CARRYB[11][27] ), .S(\SUMB[11][27] ) );
  FA_X1 S2_11_28 ( .A(\ab[11][28] ), .B(\CARRYB[10][28] ), .CI(\SUMB[10][29] ), 
        .CO(\CARRYB[11][28] ), .S(\SUMB[11][28] ) );
  FA_X1 S2_11_29 ( .A(\ab[11][29] ), .B(\CARRYB[10][29] ), .CI(\SUMB[10][30] ), 
        .CO(\CARRYB[11][29] ), .S(\SUMB[11][29] ) );
  FA_X1 S3_11_30 ( .A(\ab[11][30] ), .B(\CARRYB[10][30] ), .CI(\ab[10][31] ), 
        .CO(\CARRYB[11][30] ), .S(\SUMB[11][30] ) );
  FA_X1 S1_10_0 ( .A(\ab[10][0] ), .B(\CARRYB[9][0] ), .CI(\SUMB[9][1] ), .CO(
        \CARRYB[10][0] ), .S(\A1[8] ) );
  FA_X1 S2_10_1 ( .A(\ab[10][1] ), .B(\CARRYB[9][1] ), .CI(\SUMB[9][2] ), .CO(
        \CARRYB[10][1] ), .S(\SUMB[10][1] ) );
  FA_X1 S2_10_2 ( .A(\ab[10][2] ), .B(\CARRYB[9][2] ), .CI(\SUMB[9][3] ), .CO(
        \CARRYB[10][2] ), .S(\SUMB[10][2] ) );
  FA_X1 S2_10_3 ( .A(\ab[10][3] ), .B(\CARRYB[9][3] ), .CI(\SUMB[9][4] ), .CO(
        \CARRYB[10][3] ), .S(\SUMB[10][3] ) );
  FA_X1 S2_10_4 ( .A(\ab[10][4] ), .B(\CARRYB[9][4] ), .CI(\SUMB[9][5] ), .CO(
        \CARRYB[10][4] ), .S(\SUMB[10][4] ) );
  FA_X1 S2_10_5 ( .A(\ab[10][5] ), .B(\CARRYB[9][5] ), .CI(\SUMB[9][6] ), .CO(
        \CARRYB[10][5] ), .S(\SUMB[10][5] ) );
  FA_X1 S2_10_6 ( .A(\ab[10][6] ), .B(\CARRYB[9][6] ), .CI(\SUMB[9][7] ), .CO(
        \CARRYB[10][6] ), .S(\SUMB[10][6] ) );
  FA_X1 S2_10_7 ( .A(\ab[10][7] ), .B(\CARRYB[9][7] ), .CI(\SUMB[9][8] ), .CO(
        \CARRYB[10][7] ), .S(\SUMB[10][7] ) );
  FA_X1 S2_10_8 ( .A(\ab[10][8] ), .B(\CARRYB[9][8] ), .CI(\SUMB[9][9] ), .CO(
        \CARRYB[10][8] ), .S(\SUMB[10][8] ) );
  FA_X1 S2_10_9 ( .A(\ab[10][9] ), .B(\CARRYB[9][9] ), .CI(\SUMB[9][10] ), 
        .CO(\CARRYB[10][9] ), .S(\SUMB[10][9] ) );
  FA_X1 S2_10_10 ( .A(\ab[10][10] ), .B(\CARRYB[9][10] ), .CI(\SUMB[9][11] ), 
        .CO(\CARRYB[10][10] ), .S(\SUMB[10][10] ) );
  FA_X1 S2_10_11 ( .A(\ab[10][11] ), .B(\CARRYB[9][11] ), .CI(\SUMB[9][12] ), 
        .CO(\CARRYB[10][11] ), .S(\SUMB[10][11] ) );
  FA_X1 S2_10_12 ( .A(\ab[10][12] ), .B(\CARRYB[9][12] ), .CI(\SUMB[9][13] ), 
        .CO(\CARRYB[10][12] ), .S(\SUMB[10][12] ) );
  FA_X1 S2_10_13 ( .A(\ab[10][13] ), .B(\CARRYB[9][13] ), .CI(\SUMB[9][14] ), 
        .CO(\CARRYB[10][13] ), .S(\SUMB[10][13] ) );
  FA_X1 S2_10_14 ( .A(\ab[10][14] ), .B(\CARRYB[9][14] ), .CI(\SUMB[9][15] ), 
        .CO(\CARRYB[10][14] ), .S(\SUMB[10][14] ) );
  FA_X1 S2_10_15 ( .A(\ab[10][15] ), .B(\CARRYB[9][15] ), .CI(\SUMB[9][16] ), 
        .CO(\CARRYB[10][15] ), .S(\SUMB[10][15] ) );
  FA_X1 S2_10_16 ( .A(\ab[10][16] ), .B(\CARRYB[9][16] ), .CI(\SUMB[9][17] ), 
        .CO(\CARRYB[10][16] ), .S(\SUMB[10][16] ) );
  FA_X1 S2_10_17 ( .A(\ab[10][17] ), .B(\CARRYB[9][17] ), .CI(\SUMB[9][18] ), 
        .CO(\CARRYB[10][17] ), .S(\SUMB[10][17] ) );
  FA_X1 S2_10_18 ( .A(\ab[10][18] ), .B(\CARRYB[9][18] ), .CI(\SUMB[9][19] ), 
        .CO(\CARRYB[10][18] ), .S(\SUMB[10][18] ) );
  FA_X1 S2_10_19 ( .A(\ab[10][19] ), .B(\CARRYB[9][19] ), .CI(\SUMB[9][20] ), 
        .CO(\CARRYB[10][19] ), .S(\SUMB[10][19] ) );
  FA_X1 S2_10_20 ( .A(\CARRYB[9][20] ), .B(\ab[10][20] ), .CI(\SUMB[9][21] ), 
        .CO(\CARRYB[10][20] ), .S(\SUMB[10][20] ) );
  FA_X1 S2_10_21 ( .A(\CARRYB[9][21] ), .B(\ab[10][21] ), .CI(\SUMB[9][22] ), 
        .CO(\CARRYB[10][21] ), .S(\SUMB[10][21] ) );
  FA_X1 S2_10_26 ( .A(\ab[10][26] ), .B(\CARRYB[9][26] ), .CI(\SUMB[9][27] ), 
        .CO(\CARRYB[10][26] ), .S(\SUMB[10][26] ) );
  FA_X1 S2_10_27 ( .A(\ab[10][27] ), .B(\CARRYB[9][27] ), .CI(\SUMB[9][28] ), 
        .CO(\CARRYB[10][27] ), .S(\SUMB[10][27] ) );
  FA_X1 S2_10_28 ( .A(\ab[10][28] ), .B(\CARRYB[9][28] ), .CI(\SUMB[9][29] ), 
        .CO(\CARRYB[10][28] ), .S(\SUMB[10][28] ) );
  FA_X1 S2_10_29 ( .A(\ab[10][29] ), .B(\CARRYB[9][29] ), .CI(\SUMB[9][30] ), 
        .CO(\CARRYB[10][29] ), .S(\SUMB[10][29] ) );
  FA_X1 S3_10_30 ( .A(\ab[10][30] ), .B(\CARRYB[9][30] ), .CI(\ab[9][31] ), 
        .CO(\CARRYB[10][30] ), .S(\SUMB[10][30] ) );
  FA_X1 S1_9_0 ( .A(\ab[9][0] ), .B(\CARRYB[8][0] ), .CI(\SUMB[8][1] ), .CO(
        \CARRYB[9][0] ), .S(\A1[7] ) );
  FA_X1 S2_9_1 ( .A(\ab[9][1] ), .B(\CARRYB[8][1] ), .CI(\SUMB[8][2] ), .CO(
        \CARRYB[9][1] ), .S(\SUMB[9][1] ) );
  FA_X1 S2_9_2 ( .A(\ab[9][2] ), .B(\CARRYB[8][2] ), .CI(\SUMB[8][3] ), .CO(
        \CARRYB[9][2] ), .S(\SUMB[9][2] ) );
  FA_X1 S2_9_3 ( .A(\ab[9][3] ), .B(\CARRYB[8][3] ), .CI(\SUMB[8][4] ), .CO(
        \CARRYB[9][3] ), .S(\SUMB[9][3] ) );
  FA_X1 S2_9_4 ( .A(\ab[9][4] ), .B(\CARRYB[8][4] ), .CI(\SUMB[8][5] ), .CO(
        \CARRYB[9][4] ), .S(\SUMB[9][4] ) );
  FA_X1 S2_9_5 ( .A(\ab[9][5] ), .B(\CARRYB[8][5] ), .CI(\SUMB[8][6] ), .CO(
        \CARRYB[9][5] ), .S(\SUMB[9][5] ) );
  FA_X1 S2_9_6 ( .A(\ab[9][6] ), .B(\CARRYB[8][6] ), .CI(\SUMB[8][7] ), .CO(
        \CARRYB[9][6] ), .S(\SUMB[9][6] ) );
  FA_X1 S2_9_7 ( .A(\ab[9][7] ), .B(\CARRYB[8][7] ), .CI(\SUMB[8][8] ), .CO(
        \CARRYB[9][7] ), .S(\SUMB[9][7] ) );
  FA_X1 S2_9_8 ( .A(\ab[9][8] ), .B(\CARRYB[8][8] ), .CI(\SUMB[8][9] ), .CO(
        \CARRYB[9][8] ), .S(\SUMB[9][8] ) );
  FA_X1 S2_9_9 ( .A(\ab[9][9] ), .B(\CARRYB[8][9] ), .CI(\SUMB[8][10] ), .CO(
        \CARRYB[9][9] ), .S(\SUMB[9][9] ) );
  FA_X1 S2_9_10 ( .A(\ab[9][10] ), .B(\CARRYB[8][10] ), .CI(\SUMB[8][11] ), 
        .CO(\CARRYB[9][10] ), .S(\SUMB[9][10] ) );
  FA_X1 S2_9_11 ( .A(\ab[9][11] ), .B(\CARRYB[8][11] ), .CI(\SUMB[8][12] ), 
        .CO(\CARRYB[9][11] ), .S(\SUMB[9][11] ) );
  FA_X1 S2_9_12 ( .A(\ab[9][12] ), .B(\CARRYB[8][12] ), .CI(\SUMB[8][13] ), 
        .CO(\CARRYB[9][12] ), .S(\SUMB[9][12] ) );
  FA_X1 S2_9_13 ( .A(\ab[9][13] ), .B(\CARRYB[8][13] ), .CI(\SUMB[8][14] ), 
        .CO(\CARRYB[9][13] ), .S(\SUMB[9][13] ) );
  FA_X1 S2_9_14 ( .A(\ab[9][14] ), .B(\CARRYB[8][14] ), .CI(\SUMB[8][15] ), 
        .CO(\CARRYB[9][14] ), .S(\SUMB[9][14] ) );
  FA_X1 S2_9_15 ( .A(\ab[9][15] ), .B(\CARRYB[8][15] ), .CI(\SUMB[8][16] ), 
        .CO(\CARRYB[9][15] ), .S(\SUMB[9][15] ) );
  FA_X1 S2_9_16 ( .A(\ab[9][16] ), .B(\CARRYB[8][16] ), .CI(\SUMB[8][17] ), 
        .CO(\CARRYB[9][16] ), .S(\SUMB[9][16] ) );
  FA_X1 S2_9_17 ( .A(\ab[9][17] ), .B(\CARRYB[8][17] ), .CI(\SUMB[8][18] ), 
        .CO(\CARRYB[9][17] ), .S(\SUMB[9][17] ) );
  FA_X1 S2_9_18 ( .A(\ab[9][18] ), .B(\CARRYB[8][18] ), .CI(\SUMB[8][19] ), 
        .CO(\CARRYB[9][18] ), .S(\SUMB[9][18] ) );
  FA_X1 S2_9_19 ( .A(\ab[9][19] ), .B(\CARRYB[8][19] ), .CI(\SUMB[8][20] ), 
        .CO(\CARRYB[9][19] ), .S(\SUMB[9][19] ) );
  FA_X1 S2_9_20 ( .A(\ab[9][20] ), .B(\CARRYB[8][20] ), .CI(\SUMB[8][21] ), 
        .CO(\CARRYB[9][20] ), .S(\SUMB[9][20] ) );
  FA_X1 S2_9_21 ( .A(\CARRYB[8][21] ), .B(\ab[9][21] ), .CI(\SUMB[8][22] ), 
        .CO(\CARRYB[9][21] ), .S(\SUMB[9][21] ) );
  FA_X1 S2_9_22 ( .A(\CARRYB[8][22] ), .B(\ab[9][22] ), .CI(\SUMB[8][23] ), 
        .CO(\CARRYB[9][22] ), .S(\SUMB[9][22] ) );
  FA_X1 S2_9_27 ( .A(\ab[9][27] ), .B(\CARRYB[8][27] ), .CI(\SUMB[8][28] ), 
        .CO(\CARRYB[9][27] ), .S(\SUMB[9][27] ) );
  FA_X1 S2_9_28 ( .A(\ab[9][28] ), .B(\CARRYB[8][28] ), .CI(\SUMB[8][29] ), 
        .CO(\CARRYB[9][28] ), .S(\SUMB[9][28] ) );
  FA_X1 S2_9_29 ( .A(\ab[9][29] ), .B(\CARRYB[8][29] ), .CI(\SUMB[8][30] ), 
        .CO(\CARRYB[9][29] ), .S(\SUMB[9][29] ) );
  FA_X1 S3_9_30 ( .A(\ab[9][30] ), .B(\CARRYB[8][30] ), .CI(\ab[8][31] ), .CO(
        \CARRYB[9][30] ), .S(\SUMB[9][30] ) );
  FA_X1 S1_8_0 ( .A(\ab[8][0] ), .B(\CARRYB[7][0] ), .CI(\SUMB[7][1] ), .CO(
        \CARRYB[8][0] ), .S(\A1[6] ) );
  FA_X1 S2_8_1 ( .A(\ab[8][1] ), .B(\CARRYB[7][1] ), .CI(\SUMB[7][2] ), .CO(
        \CARRYB[8][1] ), .S(\SUMB[8][1] ) );
  FA_X1 S2_8_2 ( .A(\ab[8][2] ), .B(\CARRYB[7][2] ), .CI(\SUMB[7][3] ), .CO(
        \CARRYB[8][2] ), .S(\SUMB[8][2] ) );
  FA_X1 S2_8_3 ( .A(\ab[8][3] ), .B(\CARRYB[7][3] ), .CI(\SUMB[7][4] ), .CO(
        \CARRYB[8][3] ), .S(\SUMB[8][3] ) );
  FA_X1 S2_8_4 ( .A(\ab[8][4] ), .B(\CARRYB[7][4] ), .CI(\SUMB[7][5] ), .CO(
        \CARRYB[8][4] ), .S(\SUMB[8][4] ) );
  FA_X1 S2_8_5 ( .A(\ab[8][5] ), .B(\CARRYB[7][5] ), .CI(\SUMB[7][6] ), .CO(
        \CARRYB[8][5] ), .S(\SUMB[8][5] ) );
  FA_X1 S2_8_6 ( .A(\ab[8][6] ), .B(\CARRYB[7][6] ), .CI(\SUMB[7][7] ), .CO(
        \CARRYB[8][6] ), .S(\SUMB[8][6] ) );
  FA_X1 S2_8_7 ( .A(\ab[8][7] ), .B(\CARRYB[7][7] ), .CI(\SUMB[7][8] ), .CO(
        \CARRYB[8][7] ), .S(\SUMB[8][7] ) );
  FA_X1 S2_8_8 ( .A(\ab[8][8] ), .B(\CARRYB[7][8] ), .CI(\SUMB[7][9] ), .CO(
        \CARRYB[8][8] ), .S(\SUMB[8][8] ) );
  FA_X1 S2_8_9 ( .A(\ab[8][9] ), .B(\CARRYB[7][9] ), .CI(\SUMB[7][10] ), .CO(
        \CARRYB[8][9] ), .S(\SUMB[8][9] ) );
  FA_X1 S2_8_10 ( .A(\ab[8][10] ), .B(\CARRYB[7][10] ), .CI(\SUMB[7][11] ), 
        .CO(\CARRYB[8][10] ), .S(\SUMB[8][10] ) );
  FA_X1 S2_8_11 ( .A(\ab[8][11] ), .B(\CARRYB[7][11] ), .CI(\SUMB[7][12] ), 
        .CO(\CARRYB[8][11] ), .S(\SUMB[8][11] ) );
  FA_X1 S2_8_12 ( .A(\ab[8][12] ), .B(\CARRYB[7][12] ), .CI(\SUMB[7][13] ), 
        .CO(\CARRYB[8][12] ), .S(\SUMB[8][12] ) );
  FA_X1 S2_8_13 ( .A(\ab[8][13] ), .B(\CARRYB[7][13] ), .CI(\SUMB[7][14] ), 
        .CO(\CARRYB[8][13] ), .S(\SUMB[8][13] ) );
  FA_X1 S2_8_14 ( .A(\ab[8][14] ), .B(\CARRYB[7][14] ), .CI(\SUMB[7][15] ), 
        .CO(\CARRYB[8][14] ), .S(\SUMB[8][14] ) );
  FA_X1 S2_8_15 ( .A(\ab[8][15] ), .B(\CARRYB[7][15] ), .CI(\SUMB[7][16] ), 
        .CO(\CARRYB[8][15] ), .S(\SUMB[8][15] ) );
  FA_X1 S2_8_16 ( .A(\ab[8][16] ), .B(\CARRYB[7][16] ), .CI(\SUMB[7][17] ), 
        .CO(\CARRYB[8][16] ), .S(\SUMB[8][16] ) );
  FA_X1 S2_8_17 ( .A(\ab[8][17] ), .B(\CARRYB[7][17] ), .CI(\SUMB[7][18] ), 
        .CO(\CARRYB[8][17] ), .S(\SUMB[8][17] ) );
  FA_X1 S2_8_18 ( .A(\ab[8][18] ), .B(\CARRYB[7][18] ), .CI(\SUMB[7][19] ), 
        .CO(\CARRYB[8][18] ), .S(\SUMB[8][18] ) );
  FA_X1 S2_8_19 ( .A(\ab[8][19] ), .B(\CARRYB[7][19] ), .CI(\SUMB[7][20] ), 
        .CO(\CARRYB[8][19] ), .S(\SUMB[8][19] ) );
  FA_X1 S2_8_20 ( .A(\ab[8][20] ), .B(\CARRYB[7][20] ), .CI(\SUMB[7][21] ), 
        .CO(\CARRYB[8][20] ), .S(\SUMB[8][20] ) );
  FA_X1 S2_8_21 ( .A(\CARRYB[7][21] ), .B(\ab[8][21] ), .CI(\SUMB[7][22] ), 
        .CO(\CARRYB[8][21] ), .S(\SUMB[8][21] ) );
  FA_X1 S2_8_22 ( .A(\CARRYB[7][22] ), .B(\ab[8][22] ), .CI(\SUMB[7][23] ), 
        .CO(\CARRYB[8][22] ), .S(\SUMB[8][22] ) );
  FA_X1 S2_8_23 ( .A(\ab[8][23] ), .B(\CARRYB[7][23] ), .CI(\SUMB[7][24] ), 
        .CO(\CARRYB[8][23] ), .S(\SUMB[8][23] ) );
  FA_X1 S2_8_28 ( .A(\ab[8][28] ), .B(\CARRYB[7][28] ), .CI(\SUMB[7][29] ), 
        .CO(\CARRYB[8][28] ), .S(\SUMB[8][28] ) );
  FA_X1 S2_8_29 ( .A(\ab[8][29] ), .B(\CARRYB[7][29] ), .CI(\SUMB[7][30] ), 
        .CO(\CARRYB[8][29] ), .S(\SUMB[8][29] ) );
  FA_X1 S3_8_30 ( .A(\ab[8][30] ), .B(\CARRYB[7][30] ), .CI(\ab[7][31] ), .CO(
        \CARRYB[8][30] ), .S(\SUMB[8][30] ) );
  FA_X1 S1_7_0 ( .A(\ab[7][0] ), .B(\CARRYB[6][0] ), .CI(\SUMB[6][1] ), .CO(
        \CARRYB[7][0] ), .S(\A1[5] ) );
  FA_X1 S2_7_1 ( .A(\ab[7][1] ), .B(\CARRYB[6][1] ), .CI(\SUMB[6][2] ), .CO(
        \CARRYB[7][1] ), .S(\SUMB[7][1] ) );
  FA_X1 S2_7_2 ( .A(\ab[7][2] ), .B(\CARRYB[6][2] ), .CI(\SUMB[6][3] ), .CO(
        \CARRYB[7][2] ), .S(\SUMB[7][2] ) );
  FA_X1 S2_7_3 ( .A(\ab[7][3] ), .B(\CARRYB[6][3] ), .CI(\SUMB[6][4] ), .CO(
        \CARRYB[7][3] ), .S(\SUMB[7][3] ) );
  FA_X1 S2_7_4 ( .A(\ab[7][4] ), .B(\CARRYB[6][4] ), .CI(\SUMB[6][5] ), .CO(
        \CARRYB[7][4] ), .S(\SUMB[7][4] ) );
  FA_X1 S2_7_5 ( .A(\ab[7][5] ), .B(\CARRYB[6][5] ), .CI(\SUMB[6][6] ), .CO(
        \CARRYB[7][5] ), .S(\SUMB[7][5] ) );
  FA_X1 S2_7_6 ( .A(\ab[7][6] ), .B(\CARRYB[6][6] ), .CI(\SUMB[6][7] ), .CO(
        \CARRYB[7][6] ), .S(\SUMB[7][6] ) );
  FA_X1 S2_7_7 ( .A(\ab[7][7] ), .B(\CARRYB[6][7] ), .CI(\SUMB[6][8] ), .CO(
        \CARRYB[7][7] ), .S(\SUMB[7][7] ) );
  FA_X1 S2_7_8 ( .A(\ab[7][8] ), .B(\CARRYB[6][8] ), .CI(\SUMB[6][9] ), .CO(
        \CARRYB[7][8] ), .S(\SUMB[7][8] ) );
  FA_X1 S2_7_9 ( .A(\ab[7][9] ), .B(\CARRYB[6][9] ), .CI(\SUMB[6][10] ), .CO(
        \CARRYB[7][9] ), .S(\SUMB[7][9] ) );
  FA_X1 S2_7_10 ( .A(\ab[7][10] ), .B(\CARRYB[6][10] ), .CI(\SUMB[6][11] ), 
        .CO(\CARRYB[7][10] ), .S(\SUMB[7][10] ) );
  FA_X1 S2_7_11 ( .A(\ab[7][11] ), .B(\CARRYB[6][11] ), .CI(\SUMB[6][12] ), 
        .CO(\CARRYB[7][11] ), .S(\SUMB[7][11] ) );
  FA_X1 S2_7_12 ( .A(\ab[7][12] ), .B(\CARRYB[6][12] ), .CI(\SUMB[6][13] ), 
        .CO(\CARRYB[7][12] ), .S(\SUMB[7][12] ) );
  FA_X1 S2_7_13 ( .A(\ab[7][13] ), .B(\CARRYB[6][13] ), .CI(\SUMB[6][14] ), 
        .CO(\CARRYB[7][13] ), .S(\SUMB[7][13] ) );
  FA_X1 S2_7_14 ( .A(\ab[7][14] ), .B(\CARRYB[6][14] ), .CI(\SUMB[6][15] ), 
        .CO(\CARRYB[7][14] ), .S(\SUMB[7][14] ) );
  FA_X1 S2_7_15 ( .A(\ab[7][15] ), .B(\CARRYB[6][15] ), .CI(\SUMB[6][16] ), 
        .CO(\CARRYB[7][15] ), .S(\SUMB[7][15] ) );
  FA_X1 S2_7_16 ( .A(\ab[7][16] ), .B(\CARRYB[6][16] ), .CI(\SUMB[6][17] ), 
        .CO(\CARRYB[7][16] ), .S(\SUMB[7][16] ) );
  FA_X1 S2_7_17 ( .A(\ab[7][17] ), .B(\CARRYB[6][17] ), .CI(\SUMB[6][18] ), 
        .CO(\CARRYB[7][17] ), .S(\SUMB[7][17] ) );
  FA_X1 S2_7_18 ( .A(\ab[7][18] ), .B(\CARRYB[6][18] ), .CI(\SUMB[6][19] ), 
        .CO(\CARRYB[7][18] ), .S(\SUMB[7][18] ) );
  FA_X1 S2_7_19 ( .A(\ab[7][19] ), .B(\CARRYB[6][19] ), .CI(\SUMB[6][20] ), 
        .CO(\CARRYB[7][19] ), .S(\SUMB[7][19] ) );
  FA_X1 S2_7_20 ( .A(\ab[7][20] ), .B(\CARRYB[6][20] ), .CI(\SUMB[6][21] ), 
        .CO(\CARRYB[7][20] ), .S(\SUMB[7][20] ) );
  FA_X1 S2_7_21 ( .A(\ab[7][21] ), .B(\CARRYB[6][21] ), .CI(\SUMB[6][22] ), 
        .CO(\CARRYB[7][21] ), .S(\SUMB[7][21] ) );
  FA_X1 S2_7_22 ( .A(\ab[7][22] ), .B(\CARRYB[6][22] ), .CI(\SUMB[6][23] ), 
        .CO(\CARRYB[7][22] ), .S(\SUMB[7][22] ) );
  FA_X1 S2_7_23 ( .A(\CARRYB[6][23] ), .B(\ab[7][23] ), .CI(\SUMB[6][24] ), 
        .CO(\CARRYB[7][23] ), .S(\SUMB[7][23] ) );
  FA_X1 S2_7_24 ( .A(\CARRYB[6][24] ), .B(\ab[7][24] ), .CI(\SUMB[6][25] ), 
        .CO(\CARRYB[7][24] ), .S(\SUMB[7][24] ) );
  FA_X1 S2_7_29 ( .A(\ab[7][29] ), .B(\CARRYB[6][29] ), .CI(\SUMB[6][30] ), 
        .CO(\CARRYB[7][29] ), .S(\SUMB[7][29] ) );
  FA_X1 S3_7_30 ( .A(\ab[7][30] ), .B(\CARRYB[6][30] ), .CI(\ab[6][31] ), .CO(
        \CARRYB[7][30] ), .S(\SUMB[7][30] ) );
  FA_X1 S1_6_0 ( .A(\ab[6][0] ), .B(\CARRYB[5][0] ), .CI(\SUMB[5][1] ), .CO(
        \CARRYB[6][0] ), .S(\A1[4] ) );
  FA_X1 S2_6_1 ( .A(\ab[6][1] ), .B(\CARRYB[5][1] ), .CI(\SUMB[5][2] ), .CO(
        \CARRYB[6][1] ), .S(\SUMB[6][1] ) );
  FA_X1 S2_6_2 ( .A(\ab[6][2] ), .B(\CARRYB[5][2] ), .CI(\SUMB[5][3] ), .CO(
        \CARRYB[6][2] ), .S(\SUMB[6][2] ) );
  FA_X1 S2_6_3 ( .A(\ab[6][3] ), .B(\CARRYB[5][3] ), .CI(\SUMB[5][4] ), .CO(
        \CARRYB[6][3] ), .S(\SUMB[6][3] ) );
  FA_X1 S2_6_4 ( .A(\ab[6][4] ), .B(\CARRYB[5][4] ), .CI(\SUMB[5][5] ), .CO(
        \CARRYB[6][4] ), .S(\SUMB[6][4] ) );
  FA_X1 S2_6_5 ( .A(\ab[6][5] ), .B(\CARRYB[5][5] ), .CI(\SUMB[5][6] ), .CO(
        \CARRYB[6][5] ), .S(\SUMB[6][5] ) );
  FA_X1 S2_6_6 ( .A(\ab[6][6] ), .B(\CARRYB[5][6] ), .CI(\SUMB[5][7] ), .CO(
        \CARRYB[6][6] ), .S(\SUMB[6][6] ) );
  FA_X1 S2_6_7 ( .A(\ab[6][7] ), .B(\CARRYB[5][7] ), .CI(\SUMB[5][8] ), .CO(
        \CARRYB[6][7] ), .S(\SUMB[6][7] ) );
  FA_X1 S2_6_8 ( .A(\ab[6][8] ), .B(\CARRYB[5][8] ), .CI(\SUMB[5][9] ), .CO(
        \CARRYB[6][8] ), .S(\SUMB[6][8] ) );
  FA_X1 S2_6_9 ( .A(\ab[6][9] ), .B(\CARRYB[5][9] ), .CI(\SUMB[5][10] ), .CO(
        \CARRYB[6][9] ), .S(\SUMB[6][9] ) );
  FA_X1 S2_6_10 ( .A(\ab[6][10] ), .B(\CARRYB[5][10] ), .CI(\SUMB[5][11] ), 
        .CO(\CARRYB[6][10] ), .S(\SUMB[6][10] ) );
  FA_X1 S2_6_11 ( .A(\ab[6][11] ), .B(\CARRYB[5][11] ), .CI(\SUMB[5][12] ), 
        .CO(\CARRYB[6][11] ), .S(\SUMB[6][11] ) );
  FA_X1 S2_6_12 ( .A(\ab[6][12] ), .B(\CARRYB[5][12] ), .CI(\SUMB[5][13] ), 
        .CO(\CARRYB[6][12] ), .S(\SUMB[6][12] ) );
  FA_X1 S2_6_13 ( .A(\ab[6][13] ), .B(\CARRYB[5][13] ), .CI(\SUMB[5][14] ), 
        .CO(\CARRYB[6][13] ), .S(\SUMB[6][13] ) );
  FA_X1 S2_6_14 ( .A(\ab[6][14] ), .B(\CARRYB[5][14] ), .CI(\SUMB[5][15] ), 
        .CO(\CARRYB[6][14] ), .S(\SUMB[6][14] ) );
  FA_X1 S2_6_15 ( .A(\ab[6][15] ), .B(\CARRYB[5][15] ), .CI(\SUMB[5][16] ), 
        .CO(\CARRYB[6][15] ), .S(\SUMB[6][15] ) );
  FA_X1 S2_6_16 ( .A(\ab[6][16] ), .B(\CARRYB[5][16] ), .CI(\SUMB[5][17] ), 
        .CO(\CARRYB[6][16] ), .S(\SUMB[6][16] ) );
  FA_X1 S2_6_17 ( .A(\ab[6][17] ), .B(\CARRYB[5][17] ), .CI(\SUMB[5][18] ), 
        .CO(\CARRYB[6][17] ), .S(\SUMB[6][17] ) );
  FA_X1 S2_6_18 ( .A(\ab[6][18] ), .B(\CARRYB[5][18] ), .CI(\SUMB[5][19] ), 
        .CO(\CARRYB[6][18] ), .S(\SUMB[6][18] ) );
  FA_X1 S2_6_19 ( .A(\ab[6][19] ), .B(\CARRYB[5][19] ), .CI(\SUMB[5][20] ), 
        .CO(\CARRYB[6][19] ), .S(\SUMB[6][19] ) );
  FA_X1 S2_6_20 ( .A(\ab[6][20] ), .B(\CARRYB[5][20] ), .CI(\SUMB[5][21] ), 
        .CO(\CARRYB[6][20] ), .S(\SUMB[6][20] ) );
  FA_X1 S2_6_21 ( .A(\ab[6][21] ), .B(\CARRYB[5][21] ), .CI(\SUMB[5][22] ), 
        .CO(\CARRYB[6][21] ), .S(\SUMB[6][21] ) );
  FA_X1 S2_6_22 ( .A(\ab[6][22] ), .B(\CARRYB[5][22] ), .CI(\SUMB[5][23] ), 
        .CO(\CARRYB[6][22] ), .S(\SUMB[6][22] ) );
  FA_X1 S2_6_23 ( .A(\CARRYB[5][23] ), .B(\ab[6][23] ), .CI(\SUMB[5][24] ), 
        .CO(\CARRYB[6][23] ), .S(\SUMB[6][23] ) );
  FA_X1 S2_6_24 ( .A(\ab[6][24] ), .B(\CARRYB[5][24] ), .CI(\SUMB[5][25] ), 
        .CO(\CARRYB[6][24] ), .S(\SUMB[6][24] ) );
  FA_X1 S2_6_25 ( .A(\ab[6][25] ), .B(\CARRYB[5][25] ), .CI(\SUMB[5][26] ), 
        .CO(\CARRYB[6][25] ), .S(\SUMB[6][25] ) );
  FA_X1 S2_6_29 ( .A(\ab[6][29] ), .B(\CARRYB[5][29] ), .CI(\SUMB[5][30] ), 
        .CO(\CARRYB[6][29] ), .S(\SUMB[6][29] ) );
  FA_X1 S3_6_30 ( .A(\ab[6][30] ), .B(\CARRYB[5][30] ), .CI(\ab[5][31] ), .CO(
        \CARRYB[6][30] ), .S(\SUMB[6][30] ) );
  FA_X1 S1_5_0 ( .A(\ab[5][0] ), .B(\CARRYB[4][0] ), .CI(\SUMB[4][1] ), .CO(
        \CARRYB[5][0] ), .S(\A1[3] ) );
  FA_X1 S2_5_1 ( .A(\ab[5][1] ), .B(\CARRYB[4][1] ), .CI(\SUMB[4][2] ), .CO(
        \CARRYB[5][1] ), .S(\SUMB[5][1] ) );
  FA_X1 S2_5_2 ( .A(\ab[5][2] ), .B(\CARRYB[4][2] ), .CI(\SUMB[4][3] ), .CO(
        \CARRYB[5][2] ), .S(\SUMB[5][2] ) );
  FA_X1 S2_5_3 ( .A(\ab[5][3] ), .B(\CARRYB[4][3] ), .CI(\SUMB[4][4] ), .CO(
        \CARRYB[5][3] ), .S(\SUMB[5][3] ) );
  FA_X1 S2_5_4 ( .A(\ab[5][4] ), .B(\CARRYB[4][4] ), .CI(\SUMB[4][5] ), .CO(
        \CARRYB[5][4] ), .S(\SUMB[5][4] ) );
  FA_X1 S2_5_5 ( .A(\ab[5][5] ), .B(\CARRYB[4][5] ), .CI(\SUMB[4][6] ), .CO(
        \CARRYB[5][5] ), .S(\SUMB[5][5] ) );
  FA_X1 S2_5_6 ( .A(\ab[5][6] ), .B(\CARRYB[4][6] ), .CI(\SUMB[4][7] ), .CO(
        \CARRYB[5][6] ), .S(\SUMB[5][6] ) );
  FA_X1 S2_5_7 ( .A(\ab[5][7] ), .B(\CARRYB[4][7] ), .CI(\SUMB[4][8] ), .CO(
        \CARRYB[5][7] ), .S(\SUMB[5][7] ) );
  FA_X1 S2_5_8 ( .A(\ab[5][8] ), .B(\CARRYB[4][8] ), .CI(\SUMB[4][9] ), .CO(
        \CARRYB[5][8] ), .S(\SUMB[5][8] ) );
  FA_X1 S2_5_9 ( .A(\ab[5][9] ), .B(\CARRYB[4][9] ), .CI(\SUMB[4][10] ), .CO(
        \CARRYB[5][9] ), .S(\SUMB[5][9] ) );
  FA_X1 S2_5_10 ( .A(\ab[5][10] ), .B(\CARRYB[4][10] ), .CI(\SUMB[4][11] ), 
        .CO(\CARRYB[5][10] ), .S(\SUMB[5][10] ) );
  FA_X1 S2_5_11 ( .A(\ab[5][11] ), .B(\CARRYB[4][11] ), .CI(\SUMB[4][12] ), 
        .CO(\CARRYB[5][11] ), .S(\SUMB[5][11] ) );
  FA_X1 S2_5_12 ( .A(\ab[5][12] ), .B(\CARRYB[4][12] ), .CI(\SUMB[4][13] ), 
        .CO(\CARRYB[5][12] ), .S(\SUMB[5][12] ) );
  FA_X1 S2_5_13 ( .A(\ab[5][13] ), .B(\CARRYB[4][13] ), .CI(\SUMB[4][14] ), 
        .CO(\CARRYB[5][13] ), .S(\SUMB[5][13] ) );
  FA_X1 S2_5_14 ( .A(\ab[5][14] ), .B(\CARRYB[4][14] ), .CI(\SUMB[4][15] ), 
        .CO(\CARRYB[5][14] ), .S(\SUMB[5][14] ) );
  FA_X1 S2_5_15 ( .A(\ab[5][15] ), .B(\CARRYB[4][15] ), .CI(\SUMB[4][16] ), 
        .CO(\CARRYB[5][15] ), .S(\SUMB[5][15] ) );
  FA_X1 S2_5_16 ( .A(\ab[5][16] ), .B(\CARRYB[4][16] ), .CI(\SUMB[4][17] ), 
        .CO(\CARRYB[5][16] ), .S(\SUMB[5][16] ) );
  FA_X1 S2_5_17 ( .A(\ab[5][17] ), .B(\CARRYB[4][17] ), .CI(\SUMB[4][18] ), 
        .CO(\CARRYB[5][17] ), .S(\SUMB[5][17] ) );
  FA_X1 S2_5_18 ( .A(\ab[5][18] ), .B(\CARRYB[4][18] ), .CI(\SUMB[4][19] ), 
        .CO(\CARRYB[5][18] ), .S(\SUMB[5][18] ) );
  FA_X1 S2_5_19 ( .A(\ab[5][19] ), .B(\CARRYB[4][19] ), .CI(\SUMB[4][20] ), 
        .CO(\CARRYB[5][19] ), .S(\SUMB[5][19] ) );
  FA_X1 S2_5_20 ( .A(\ab[5][20] ), .B(\CARRYB[4][20] ), .CI(\SUMB[4][21] ), 
        .CO(\CARRYB[5][20] ), .S(\SUMB[5][20] ) );
  FA_X1 S2_5_21 ( .A(\ab[5][21] ), .B(\CARRYB[4][21] ), .CI(\SUMB[4][22] ), 
        .CO(\CARRYB[5][21] ), .S(\SUMB[5][21] ) );
  FA_X1 S2_5_22 ( .A(\ab[5][22] ), .B(\CARRYB[4][22] ), .CI(\SUMB[4][23] ), 
        .CO(\CARRYB[5][22] ), .S(\SUMB[5][22] ) );
  FA_X1 S2_5_23 ( .A(\ab[5][23] ), .B(\CARRYB[4][23] ), .CI(\SUMB[4][24] ), 
        .CO(\CARRYB[5][23] ), .S(\SUMB[5][23] ) );
  FA_X1 S2_5_24 ( .A(\ab[5][24] ), .B(\CARRYB[4][24] ), .CI(\SUMB[4][25] ), 
        .CO(\CARRYB[5][24] ), .S(\SUMB[5][24] ) );
  FA_X1 S2_5_25 ( .A(\CARRYB[4][25] ), .B(\ab[5][25] ), .CI(\SUMB[4][26] ), 
        .CO(\CARRYB[5][25] ), .S(\SUMB[5][25] ) );
  FA_X1 S2_5_26 ( .A(\ab[5][26] ), .B(\CARRYB[4][26] ), .CI(\SUMB[4][27] ), 
        .CO(\CARRYB[5][26] ), .S(\SUMB[5][26] ) );
  FA_X1 S3_5_30 ( .A(\ab[5][30] ), .B(\CARRYB[4][30] ), .CI(\ab[4][31] ), .CO(
        \CARRYB[5][30] ), .S(\SUMB[5][30] ) );
  FA_X1 S1_4_0 ( .A(\ab[4][0] ), .B(\CARRYB[3][0] ), .CI(\SUMB[3][1] ), .CO(
        \CARRYB[4][0] ), .S(\A1[2] ) );
  FA_X1 S2_4_1 ( .A(\ab[4][1] ), .B(\CARRYB[3][1] ), .CI(\SUMB[3][2] ), .CO(
        \CARRYB[4][1] ), .S(\SUMB[4][1] ) );
  FA_X1 S2_4_2 ( .A(\ab[4][2] ), .B(\CARRYB[3][2] ), .CI(\SUMB[3][3] ), .CO(
        \CARRYB[4][2] ), .S(\SUMB[4][2] ) );
  FA_X1 S2_4_3 ( .A(\ab[4][3] ), .B(\CARRYB[3][3] ), .CI(\SUMB[3][4] ), .CO(
        \CARRYB[4][3] ), .S(\SUMB[4][3] ) );
  FA_X1 S2_4_4 ( .A(\ab[4][4] ), .B(\CARRYB[3][4] ), .CI(\SUMB[3][5] ), .CO(
        \CARRYB[4][4] ), .S(\SUMB[4][4] ) );
  FA_X1 S2_4_5 ( .A(\ab[4][5] ), .B(\CARRYB[3][5] ), .CI(\SUMB[3][6] ), .CO(
        \CARRYB[4][5] ), .S(\SUMB[4][5] ) );
  FA_X1 S2_4_6 ( .A(\ab[4][6] ), .B(\CARRYB[3][6] ), .CI(\SUMB[3][7] ), .CO(
        \CARRYB[4][6] ), .S(\SUMB[4][6] ) );
  FA_X1 S2_4_7 ( .A(\ab[4][7] ), .B(\CARRYB[3][7] ), .CI(\SUMB[3][8] ), .CO(
        \CARRYB[4][7] ), .S(\SUMB[4][7] ) );
  FA_X1 S2_4_8 ( .A(\ab[4][8] ), .B(\CARRYB[3][8] ), .CI(\SUMB[3][9] ), .CO(
        \CARRYB[4][8] ), .S(\SUMB[4][8] ) );
  FA_X1 S2_4_9 ( .A(\ab[4][9] ), .B(\CARRYB[3][9] ), .CI(\SUMB[3][10] ), .CO(
        \CARRYB[4][9] ), .S(\SUMB[4][9] ) );
  FA_X1 S2_4_10 ( .A(\ab[4][10] ), .B(\CARRYB[3][10] ), .CI(\SUMB[3][11] ), 
        .CO(\CARRYB[4][10] ), .S(\SUMB[4][10] ) );
  FA_X1 S2_4_11 ( .A(\ab[4][11] ), .B(\CARRYB[3][11] ), .CI(\SUMB[3][12] ), 
        .CO(\CARRYB[4][11] ), .S(\SUMB[4][11] ) );
  FA_X1 S2_4_12 ( .A(\ab[4][12] ), .B(\CARRYB[3][12] ), .CI(\SUMB[3][13] ), 
        .CO(\CARRYB[4][12] ), .S(\SUMB[4][12] ) );
  FA_X1 S2_4_13 ( .A(\ab[4][13] ), .B(\CARRYB[3][13] ), .CI(\SUMB[3][14] ), 
        .CO(\CARRYB[4][13] ), .S(\SUMB[4][13] ) );
  FA_X1 S2_4_14 ( .A(\ab[4][14] ), .B(\CARRYB[3][14] ), .CI(\SUMB[3][15] ), 
        .CO(\CARRYB[4][14] ), .S(\SUMB[4][14] ) );
  FA_X1 S2_4_15 ( .A(\ab[4][15] ), .B(\CARRYB[3][15] ), .CI(\SUMB[3][16] ), 
        .CO(\CARRYB[4][15] ), .S(\SUMB[4][15] ) );
  FA_X1 S2_4_16 ( .A(\ab[4][16] ), .B(\CARRYB[3][16] ), .CI(\SUMB[3][17] ), 
        .CO(\CARRYB[4][16] ), .S(\SUMB[4][16] ) );
  FA_X1 S2_4_17 ( .A(\ab[4][17] ), .B(\CARRYB[3][17] ), .CI(\SUMB[3][18] ), 
        .CO(\CARRYB[4][17] ), .S(\SUMB[4][17] ) );
  FA_X1 S2_4_18 ( .A(\ab[4][18] ), .B(\CARRYB[3][18] ), .CI(\SUMB[3][19] ), 
        .CO(\CARRYB[4][18] ), .S(\SUMB[4][18] ) );
  FA_X1 S2_4_19 ( .A(\ab[4][19] ), .B(\CARRYB[3][19] ), .CI(\SUMB[3][20] ), 
        .CO(\CARRYB[4][19] ), .S(\SUMB[4][19] ) );
  FA_X1 S2_4_20 ( .A(\ab[4][20] ), .B(\CARRYB[3][20] ), .CI(\SUMB[3][21] ), 
        .CO(\CARRYB[4][20] ), .S(\SUMB[4][20] ) );
  FA_X1 S2_4_21 ( .A(\ab[4][21] ), .B(\CARRYB[3][21] ), .CI(\SUMB[3][22] ), 
        .CO(\CARRYB[4][21] ), .S(\SUMB[4][21] ) );
  FA_X1 S2_4_22 ( .A(\ab[4][22] ), .B(\CARRYB[3][22] ), .CI(\SUMB[3][23] ), 
        .CO(\CARRYB[4][22] ), .S(\SUMB[4][22] ) );
  FA_X1 S2_4_23 ( .A(\ab[4][23] ), .B(\CARRYB[3][23] ), .CI(\SUMB[3][24] ), 
        .CO(\CARRYB[4][23] ), .S(\SUMB[4][23] ) );
  FA_X1 S2_4_24 ( .A(\ab[4][24] ), .B(\CARRYB[3][24] ), .CI(\SUMB[3][25] ), 
        .CO(\CARRYB[4][24] ), .S(\SUMB[4][24] ) );
  FA_X1 S2_4_25 ( .A(\CARRYB[3][25] ), .B(\ab[4][25] ), .CI(\SUMB[3][26] ), 
        .CO(\CARRYB[4][25] ), .S(\SUMB[4][25] ) );
  FA_X1 S2_4_26 ( .A(\ab[4][26] ), .B(\CARRYB[3][26] ), .CI(\SUMB[3][27] ), 
        .CO(\CARRYB[4][26] ), .S(\SUMB[4][26] ) );
  FA_X1 S2_4_27 ( .A(\ab[4][27] ), .B(\CARRYB[3][27] ), .CI(\SUMB[3][28] ), 
        .CO(\CARRYB[4][27] ), .S(\SUMB[4][27] ) );
  FA_X1 S3_4_30 ( .A(\ab[4][30] ), .B(\CARRYB[3][30] ), .CI(\ab[3][31] ), .CO(
        \CARRYB[4][30] ), .S(\SUMB[4][30] ) );
  FA_X1 S1_3_0 ( .A(\ab[3][0] ), .B(\CARRYB[2][0] ), .CI(\SUMB[2][1] ), .CO(
        \CARRYB[3][0] ), .S(\A1[1] ) );
  FA_X1 S2_3_1 ( .A(\ab[3][1] ), .B(\CARRYB[2][1] ), .CI(\SUMB[2][2] ), .CO(
        \CARRYB[3][1] ), .S(\SUMB[3][1] ) );
  FA_X1 S2_3_2 ( .A(\ab[3][2] ), .B(\CARRYB[2][2] ), .CI(\SUMB[2][3] ), .CO(
        \CARRYB[3][2] ), .S(\SUMB[3][2] ) );
  FA_X1 S2_3_3 ( .A(\ab[3][3] ), .B(\CARRYB[2][3] ), .CI(\SUMB[2][4] ), .CO(
        \CARRYB[3][3] ), .S(\SUMB[3][3] ) );
  FA_X1 S2_3_4 ( .A(\ab[3][4] ), .B(\CARRYB[2][4] ), .CI(\SUMB[2][5] ), .CO(
        \CARRYB[3][4] ), .S(\SUMB[3][4] ) );
  FA_X1 S2_3_5 ( .A(\ab[3][5] ), .B(\CARRYB[2][5] ), .CI(\SUMB[2][6] ), .CO(
        \CARRYB[3][5] ), .S(\SUMB[3][5] ) );
  FA_X1 S2_3_6 ( .A(\ab[3][6] ), .B(\CARRYB[2][6] ), .CI(\SUMB[2][7] ), .CO(
        \CARRYB[3][6] ), .S(\SUMB[3][6] ) );
  FA_X1 S2_3_7 ( .A(\ab[3][7] ), .B(\CARRYB[2][7] ), .CI(\SUMB[2][8] ), .CO(
        \CARRYB[3][7] ), .S(\SUMB[3][7] ) );
  FA_X1 S2_3_8 ( .A(\ab[3][8] ), .B(\CARRYB[2][8] ), .CI(\SUMB[2][9] ), .CO(
        \CARRYB[3][8] ), .S(\SUMB[3][8] ) );
  FA_X1 S2_3_9 ( .A(\ab[3][9] ), .B(\CARRYB[2][9] ), .CI(\SUMB[2][10] ), .CO(
        \CARRYB[3][9] ), .S(\SUMB[3][9] ) );
  FA_X1 S2_3_10 ( .A(\ab[3][10] ), .B(\CARRYB[2][10] ), .CI(\SUMB[2][11] ), 
        .CO(\CARRYB[3][10] ), .S(\SUMB[3][10] ) );
  FA_X1 S2_3_11 ( .A(\ab[3][11] ), .B(\CARRYB[2][11] ), .CI(\SUMB[2][12] ), 
        .CO(\CARRYB[3][11] ), .S(\SUMB[3][11] ) );
  FA_X1 S2_3_12 ( .A(\ab[3][12] ), .B(\CARRYB[2][12] ), .CI(\SUMB[2][13] ), 
        .CO(\CARRYB[3][12] ), .S(\SUMB[3][12] ) );
  FA_X1 S2_3_13 ( .A(\ab[3][13] ), .B(\CARRYB[2][13] ), .CI(\SUMB[2][14] ), 
        .CO(\CARRYB[3][13] ), .S(\SUMB[3][13] ) );
  FA_X1 S2_3_14 ( .A(\ab[3][14] ), .B(\CARRYB[2][14] ), .CI(\SUMB[2][15] ), 
        .CO(\CARRYB[3][14] ), .S(\SUMB[3][14] ) );
  FA_X1 S2_3_15 ( .A(\ab[3][15] ), .B(\CARRYB[2][15] ), .CI(\SUMB[2][16] ), 
        .CO(\CARRYB[3][15] ), .S(\SUMB[3][15] ) );
  FA_X1 S2_3_16 ( .A(\ab[3][16] ), .B(\CARRYB[2][16] ), .CI(\SUMB[2][17] ), 
        .CO(\CARRYB[3][16] ), .S(\SUMB[3][16] ) );
  FA_X1 S2_3_17 ( .A(\ab[3][17] ), .B(\CARRYB[2][17] ), .CI(\SUMB[2][18] ), 
        .CO(\CARRYB[3][17] ), .S(\SUMB[3][17] ) );
  FA_X1 S2_3_18 ( .A(\ab[3][18] ), .B(\CARRYB[2][18] ), .CI(\SUMB[2][19] ), 
        .CO(\CARRYB[3][18] ), .S(\SUMB[3][18] ) );
  FA_X1 S2_3_19 ( .A(\ab[3][19] ), .B(\CARRYB[2][19] ), .CI(\SUMB[2][20] ), 
        .CO(\CARRYB[3][19] ), .S(\SUMB[3][19] ) );
  FA_X1 S2_3_20 ( .A(\ab[3][20] ), .B(\CARRYB[2][20] ), .CI(\SUMB[2][21] ), 
        .CO(\CARRYB[3][20] ), .S(\SUMB[3][20] ) );
  FA_X1 S2_3_21 ( .A(\ab[3][21] ), .B(\CARRYB[2][21] ), .CI(\SUMB[2][22] ), 
        .CO(\CARRYB[3][21] ), .S(\SUMB[3][21] ) );
  FA_X1 S2_3_22 ( .A(\ab[3][22] ), .B(\CARRYB[2][22] ), .CI(\SUMB[2][23] ), 
        .CO(\CARRYB[3][22] ), .S(\SUMB[3][22] ) );
  FA_X1 S2_3_23 ( .A(\ab[3][23] ), .B(\CARRYB[2][23] ), .CI(\SUMB[2][24] ), 
        .CO(\CARRYB[3][23] ), .S(\SUMB[3][23] ) );
  FA_X1 S2_3_24 ( .A(\CARRYB[2][24] ), .B(\ab[3][24] ), .CI(\SUMB[2][25] ), 
        .CO(\CARRYB[3][24] ), .S(\SUMB[3][24] ) );
  FA_X1 S2_3_25 ( .A(\SUMB[2][26] ), .B(\ab[3][25] ), .CI(\CARRYB[2][25] ), 
        .CO(\CARRYB[3][25] ), .S(\SUMB[3][25] ) );
  FA_X1 S2_3_26 ( .A(\ab[3][26] ), .B(\CARRYB[2][26] ), .CI(\SUMB[2][27] ), 
        .CO(\CARRYB[3][26] ), .S(\SUMB[3][26] ) );
  FA_X1 S2_3_27 ( .A(\CARRYB[2][27] ), .B(\ab[3][27] ), .CI(\SUMB[2][28] ), 
        .CO(\CARRYB[3][27] ), .S(\SUMB[3][27] ) );
  FA_X1 S2_3_28 ( .A(\ab[3][28] ), .B(\CARRYB[2][28] ), .CI(\SUMB[2][29] ), 
        .CO(\CARRYB[3][28] ), .S(\SUMB[3][28] ) );
  FA_X1 S1_2_0 ( .A(\ab[2][0] ), .B(\CARRYB[1][0] ), .CI(\SUMB[1][1] ), .CO(
        \CARRYB[2][0] ), .S(\A1[0] ) );
  FA_X1 S2_2_1 ( .A(\ab[2][1] ), .B(\CARRYB[1][1] ), .CI(\SUMB[1][2] ), .CO(
        \CARRYB[2][1] ), .S(\SUMB[2][1] ) );
  FA_X1 S2_2_2 ( .A(\ab[2][2] ), .B(\CARRYB[1][2] ), .CI(\SUMB[1][3] ), .CO(
        \CARRYB[2][2] ), .S(\SUMB[2][2] ) );
  FA_X1 S2_2_3 ( .A(\ab[2][3] ), .B(\CARRYB[1][3] ), .CI(\SUMB[1][4] ), .CO(
        \CARRYB[2][3] ), .S(\SUMB[2][3] ) );
  FA_X1 S2_2_4 ( .A(\ab[2][4] ), .B(\CARRYB[1][4] ), .CI(\SUMB[1][5] ), .CO(
        \CARRYB[2][4] ), .S(\SUMB[2][4] ) );
  FA_X1 S2_2_5 ( .A(\ab[2][5] ), .B(\CARRYB[1][5] ), .CI(\SUMB[1][6] ), .CO(
        \CARRYB[2][5] ), .S(\SUMB[2][5] ) );
  FA_X1 S2_2_6 ( .A(\ab[2][6] ), .B(\CARRYB[1][6] ), .CI(\SUMB[1][7] ), .CO(
        \CARRYB[2][6] ), .S(\SUMB[2][6] ) );
  FA_X1 S2_2_7 ( .A(\ab[2][7] ), .B(\CARRYB[1][7] ), .CI(\SUMB[1][8] ), .CO(
        \CARRYB[2][7] ), .S(\SUMB[2][7] ) );
  FA_X1 S2_2_8 ( .A(\ab[2][8] ), .B(\CARRYB[1][8] ), .CI(\SUMB[1][9] ), .CO(
        \CARRYB[2][8] ), .S(\SUMB[2][8] ) );
  FA_X1 S2_2_9 ( .A(\ab[2][9] ), .B(\CARRYB[1][9] ), .CI(\SUMB[1][10] ), .CO(
        \CARRYB[2][9] ), .S(\SUMB[2][9] ) );
  FA_X1 S2_2_10 ( .A(\ab[2][10] ), .B(\CARRYB[1][10] ), .CI(\SUMB[1][11] ), 
        .CO(\CARRYB[2][10] ), .S(\SUMB[2][10] ) );
  FA_X1 S2_2_11 ( .A(\ab[2][11] ), .B(\CARRYB[1][11] ), .CI(\SUMB[1][12] ), 
        .CO(\CARRYB[2][11] ), .S(\SUMB[2][11] ) );
  FA_X1 S2_2_12 ( .A(\ab[2][12] ), .B(\CARRYB[1][12] ), .CI(\SUMB[1][13] ), 
        .CO(\CARRYB[2][12] ), .S(\SUMB[2][12] ) );
  FA_X1 S2_2_13 ( .A(\ab[2][13] ), .B(\CARRYB[1][13] ), .CI(\SUMB[1][14] ), 
        .CO(\CARRYB[2][13] ), .S(\SUMB[2][13] ) );
  FA_X1 S2_2_14 ( .A(\ab[2][14] ), .B(\CARRYB[1][14] ), .CI(\SUMB[1][15] ), 
        .CO(\CARRYB[2][14] ), .S(\SUMB[2][14] ) );
  FA_X1 S2_2_15 ( .A(\ab[2][15] ), .B(\CARRYB[1][15] ), .CI(\SUMB[1][16] ), 
        .CO(\CARRYB[2][15] ), .S(\SUMB[2][15] ) );
  FA_X1 S2_2_16 ( .A(\ab[2][16] ), .B(\CARRYB[1][16] ), .CI(\SUMB[1][17] ), 
        .CO(\CARRYB[2][16] ), .S(\SUMB[2][16] ) );
  FA_X1 S2_2_17 ( .A(\ab[2][17] ), .B(\CARRYB[1][17] ), .CI(\SUMB[1][18] ), 
        .CO(\CARRYB[2][17] ), .S(\SUMB[2][17] ) );
  FA_X1 S2_2_18 ( .A(\ab[2][18] ), .B(\CARRYB[1][18] ), .CI(\SUMB[1][19] ), 
        .CO(\CARRYB[2][18] ), .S(\SUMB[2][18] ) );
  FA_X1 S2_2_19 ( .A(\ab[2][19] ), .B(\CARRYB[1][19] ), .CI(\SUMB[1][20] ), 
        .CO(\CARRYB[2][19] ), .S(\SUMB[2][19] ) );
  FA_X1 S2_2_20 ( .A(\ab[2][20] ), .B(\CARRYB[1][20] ), .CI(\SUMB[1][21] ), 
        .CO(\CARRYB[2][20] ), .S(\SUMB[2][20] ) );
  FA_X1 S2_2_21 ( .A(\ab[2][21] ), .B(\CARRYB[1][21] ), .CI(\SUMB[1][22] ), 
        .CO(\CARRYB[2][21] ), .S(\SUMB[2][21] ) );
  FA_X1 S2_2_22 ( .A(\ab[2][22] ), .B(\CARRYB[1][22] ), .CI(\SUMB[1][23] ), 
        .CO(\CARRYB[2][22] ), .S(\SUMB[2][22] ) );
  FA_X1 S2_2_23 ( .A(\ab[2][23] ), .B(\CARRYB[1][23] ), .CI(\SUMB[1][24] ), 
        .CO(\CARRYB[2][23] ), .S(\SUMB[2][23] ) );
  FA_X1 S2_2_24 ( .A(\ab[2][24] ), .B(\CARRYB[1][24] ), .CI(\SUMB[1][25] ), 
        .CO(\CARRYB[2][24] ), .S(\SUMB[2][24] ) );
  FA_X1 S2_2_25 ( .A(\CARRYB[1][25] ), .B(\ab[2][25] ), .CI(\SUMB[1][26] ), 
        .CO(\CARRYB[2][25] ), .S(\SUMB[2][25] ) );
  FA_X1 S2_2_26 ( .A(\ab[2][26] ), .B(\CARRYB[1][26] ), .CI(\SUMB[1][27] ), 
        .CO(\CARRYB[2][26] ), .S(\SUMB[2][26] ) );
  FA_X1 S2_2_27 ( .A(\ab[2][27] ), .B(\CARRYB[1][27] ), .CI(\SUMB[1][28] ), 
        .CO(\CARRYB[2][27] ), .S(\SUMB[2][27] ) );
  FA_X1 S2_2_28 ( .A(\ab[2][28] ), .B(\CARRYB[1][28] ), .CI(\SUMB[1][29] ), 
        .CO(\CARRYB[2][28] ), .S(\SUMB[2][28] ) );
  FA_X1 S2_2_29 ( .A(\CARRYB[1][29] ), .B(\ab[2][29] ), .CI(\SUMB[1][30] ), 
        .CO(\CARRYB[2][29] ), .S(\SUMB[2][29] ) );
  XOR2_X1 U67 ( .A(\CARRYB[31][10] ), .B(\SUMB[31][11] ), .Z(\A1[40] ) );
  XOR2_X1 U69 ( .A(\CARRYB[31][11] ), .B(\SUMB[31][12] ), .Z(\A1[41] ) );
  XOR2_X1 U71 ( .A(\CARRYB[31][13] ), .B(\SUMB[31][14] ), .Z(\A1[43] ) );
  XOR2_X1 U73 ( .A(\CARRYB[31][12] ), .B(\SUMB[31][13] ), .Z(\A1[42] ) );
  XOR2_X1 U76 ( .A(\CARRYB[31][0] ), .B(\SUMB[31][1] ), .Z(\A1[30] ) );
  XOR2_X1 U78 ( .A(\ab[1][0] ), .B(\ab[0][1] ), .Z(PRODUCT[1]) );
  XOR2_X1 U80 ( .A(\CARRYB[31][1] ), .B(\SUMB[31][2] ), .Z(\A1[31] ) );
  XOR2_X1 U82 ( .A(\ab[1][1] ), .B(\ab[0][2] ), .Z(\SUMB[1][1] ) );
  XOR2_X1 U88 ( .A(\ab[1][3] ), .B(\ab[0][4] ), .Z(\SUMB[1][3] ) );
  XOR2_X1 U90 ( .A(\ab[1][2] ), .B(\ab[0][3] ), .Z(\SUMB[1][2] ) );
  XOR2_X1 U92 ( .A(\CARRYB[31][4] ), .B(\SUMB[31][5] ), .Z(\A1[34] ) );
  XOR2_X1 U94 ( .A(\ab[1][4] ), .B(\ab[0][5] ), .Z(\SUMB[1][4] ) );
  XOR2_X1 U96 ( .A(\CARRYB[31][5] ), .B(\SUMB[31][6] ), .Z(\A1[35] ) );
  XOR2_X1 U98 ( .A(\ab[1][5] ), .B(\ab[0][6] ), .Z(\SUMB[1][5] ) );
  XOR2_X1 U100 ( .A(\CARRYB[31][6] ), .B(\SUMB[31][7] ), .Z(\A1[36] ) );
  XOR2_X1 U102 ( .A(\ab[1][6] ), .B(\ab[0][7] ), .Z(\SUMB[1][6] ) );
  XOR2_X1 U104 ( .A(\CARRYB[31][7] ), .B(\SUMB[31][8] ), .Z(\A1[37] ) );
  XOR2_X1 U106 ( .A(\ab[1][7] ), .B(\ab[0][8] ), .Z(\SUMB[1][7] ) );
  XOR2_X1 U108 ( .A(\CARRYB[31][9] ), .B(\SUMB[31][10] ), .Z(\A1[39] ) );
  XOR2_X1 U110 ( .A(\CARRYB[31][8] ), .B(\SUMB[31][9] ), .Z(\A1[38] ) );
  XOR2_X1 U112 ( .A(\ab[1][13] ), .B(\ab[0][14] ), .Z(\SUMB[1][13] ) );
  XOR2_X1 U114 ( .A(\ab[1][12] ), .B(\ab[0][13] ), .Z(\SUMB[1][12] ) );
  XOR2_X1 U116 ( .A(\ab[1][11] ), .B(\ab[0][12] ), .Z(\SUMB[1][11] ) );
  XOR2_X1 U118 ( .A(\ab[1][10] ), .B(\ab[0][11] ), .Z(\SUMB[1][10] ) );
  XOR2_X1 U120 ( .A(\ab[1][9] ), .B(\ab[0][10] ), .Z(\SUMB[1][9] ) );
  XOR2_X1 U122 ( .A(\ab[1][8] ), .B(\ab[0][9] ), .Z(\SUMB[1][8] ) );
  XOR2_X1 U124 ( .A(\CARRYB[31][15] ), .B(\SUMB[31][16] ), .Z(\A1[45] ) );
  XOR2_X1 U126 ( .A(\CARRYB[31][14] ), .B(\SUMB[31][15] ), .Z(\A1[44] ) );
  XOR2_X1 U128 ( .A(\ab[1][15] ), .B(\ab[0][16] ), .Z(\SUMB[1][15] ) );
  XOR2_X1 U130 ( .A(\ab[1][14] ), .B(\ab[0][15] ), .Z(\SUMB[1][14] ) );
  XOR2_X1 U132 ( .A(\CARRYB[31][16] ), .B(\SUMB[31][17] ), .Z(\A1[46] ) );
  XOR2_X1 U134 ( .A(\ab[1][16] ), .B(\ab[0][17] ), .Z(\SUMB[1][16] ) );
  XOR2_X1 U136 ( .A(\CARRYB[31][17] ), .B(\SUMB[31][18] ), .Z(\A1[47] ) );
  XOR2_X1 U138 ( .A(\ab[1][17] ), .B(\ab[0][18] ), .Z(\SUMB[1][17] ) );
  XOR2_X1 U140 ( .A(\CARRYB[31][18] ), .B(\SUMB[31][19] ), .Z(\A1[48] ) );
  XOR2_X1 U142 ( .A(\ab[1][18] ), .B(\ab[0][19] ), .Z(\SUMB[1][18] ) );
  XOR2_X1 U144 ( .A(\CARRYB[31][19] ), .B(\SUMB[31][20] ), .Z(\A1[49] ) );
  XOR2_X1 U146 ( .A(\ab[1][19] ), .B(\ab[0][20] ), .Z(\SUMB[1][19] ) );
  XOR2_X1 U148 ( .A(\CARRYB[31][20] ), .B(\SUMB[31][21] ), .Z(\A1[50] ) );
  XOR2_X1 U150 ( .A(\ab[1][20] ), .B(\ab[0][21] ), .Z(\SUMB[1][20] ) );
  XOR2_X1 U152 ( .A(\CARRYB[31][21] ), .B(\SUMB[31][22] ), .Z(\A1[51] ) );
  XOR2_X1 U154 ( .A(\ab[1][21] ), .B(\ab[0][22] ), .Z(\SUMB[1][21] ) );
  XOR2_X1 U156 ( .A(\CARRYB[31][22] ), .B(\SUMB[31][23] ), .Z(\A1[52] ) );
  XOR2_X1 U158 ( .A(\ab[1][22] ), .B(\ab[0][23] ), .Z(\SUMB[1][22] ) );
  XOR2_X1 U160 ( .A(\CARRYB[31][23] ), .B(\SUMB[31][24] ), .Z(\A1[53] ) );
  XOR2_X1 U162 ( .A(\ab[1][23] ), .B(\ab[0][24] ), .Z(\SUMB[1][23] ) );
  XOR2_X1 U164 ( .A(\CARRYB[31][24] ), .B(\SUMB[31][25] ), .Z(\A1[54] ) );
  XOR2_X1 U168 ( .A(\CARRYB[31][25] ), .B(\SUMB[31][26] ), .Z(\A1[55] ) );
  XOR2_X1 U172 ( .A(\CARRYB[31][26] ), .B(\SUMB[31][27] ), .Z(\A1[56] ) );
  XOR2_X1 U174 ( .A(\ab[1][26] ), .B(\ab[0][27] ), .Z(\SUMB[1][26] ) );
  XOR2_X1 U176 ( .A(\CARRYB[31][27] ), .B(\SUMB[31][28] ), .Z(\A1[57] ) );
  XOR2_X1 U180 ( .A(\CARRYB[31][28] ), .B(\SUMB[31][29] ), .Z(\A1[58] ) );
  XOR2_X1 U182 ( .A(\ab[1][28] ), .B(\ab[0][29] ), .Z(\SUMB[1][28] ) );
  XOR2_X1 U184 ( .A(\CARRYB[31][30] ), .B(\SUMB[31][31] ), .Z(\A1[60] ) );
  XOR2_X1 U187 ( .A(\CARRYB[31][29] ), .B(\SUMB[31][30] ), .Z(\A1[59] ) );
  Multiplier_NBIT_DATA32_DW01_add_0 FS_1 ( .A({1'b0, \A1[60] , \A1[59] , 
        \A1[58] , \A1[57] , \A1[56] , \A1[55] , \A1[54] , \A1[53] , \A1[52] , 
        \A1[51] , \A1[50] , \A1[49] , \A1[48] , \A1[47] , \A1[46] , \A1[45] , 
        \A1[44] , \A1[43] , \A1[42] , \A1[41] , \A1[40] , \A1[39] , \A1[38] , 
        \A1[37] , \A1[36] , \A1[35] , \A1[34] , \A1[33] , \A1[32] , \A1[31] , 
        \A1[30] , \A1[29] , \A1[28] , \A1[27] , \A1[26] , \A1[25] , \A1[24] , 
        \A1[23] , \A1[22] , \A1[21] , \A1[20] , \A1[19] , \A1[18] , \A1[17] , 
        \A1[16] , \A1[15] , \A1[14] , \A1[13] , \A1[12] , \A1[11] , \A1[10] , 
        \A1[9] , \A1[8] , \A1[7] , \A1[6] , \A1[5] , \A1[4] , \A1[3] , \A1[2] , 
        \A1[1] , \A1[0] }), .B({\A2[61] , \A2[60] , \A2[59] , \A2[58] , 
        \A2[57] , \A2[56] , \A2[55] , \A2[54] , \A2[53] , \A2[52] , \A2[51] , 
        \A2[50] , \A2[49] , \A2[48] , \A2[47] , \A2[46] , \A2[45] , \A2[44] , 
        \A2[43] , \A2[42] , \A2[41] , \A2[40] , \A2[39] , \A2[38] , \A2[37] , 
        \A2[36] , \A2[35] , \A2[34] , \A2[33] , \A2[32] , \A2[31] , 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM(PRODUCT[63:2]) );
  XOR2_X1 U86 ( .A(\SUMB[31][3] ), .B(\CARRYB[31][2] ), .Z(\A1[32] ) );
  XOR2_X1 U84 ( .A(\SUMB[31][4] ), .B(\CARRYB[31][3] ), .Z(\A1[33] ) );
  FA_X1 S2_18_14 ( .A(\ab[18][14] ), .B(\CARRYB[17][14] ), .CI(\SUMB[17][15] ), 
        .CO(\CARRYB[18][14] ), .S(\SUMB[18][14] ) );
  FA_X1 S4_3 ( .A(\CARRYB[30][3] ), .B(\ab[31][3] ), .CI(\SUMB[30][4] ), .CO(
        \CARRYB[31][3] ), .S(\SUMB[31][3] ) );
  FA_X1 S4_4 ( .A(\CARRYB[30][4] ), .B(\ab[31][4] ), .CI(\SUMB[30][5] ), .CO(
        \CARRYB[31][4] ), .S(\SUMB[31][4] ) );
  FA_X1 S2_30_4 ( .A(\CARRYB[29][4] ), .B(\ab[30][4] ), .CI(\SUMB[29][5] ), 
        .CO(\CARRYB[30][4] ), .S(\SUMB[30][4] ) );
  FA_X1 S2_30_5 ( .A(\CARRYB[29][5] ), .B(\ab[30][5] ), .CI(\SUMB[29][6] ), 
        .CO(\CARRYB[30][5] ), .S(\SUMB[30][5] ) );
  FA_X1 S2_29_5 ( .A(\CARRYB[28][5] ), .B(\ab[29][5] ), .CI(\SUMB[28][6] ), 
        .CO(\CARRYB[29][5] ), .S(\SUMB[29][5] ) );
  FA_X1 S2_29_6 ( .A(\CARRYB[28][6] ), .B(\ab[29][6] ), .CI(\SUMB[28][7] ), 
        .CO(\CARRYB[29][6] ), .S(\SUMB[29][6] ) );
  FA_X1 S2_28_6 ( .A(\CARRYB[27][6] ), .B(\ab[28][6] ), .CI(\SUMB[27][7] ), 
        .CO(\CARRYB[28][6] ), .S(\SUMB[28][6] ) );
  FA_X1 S2_28_7 ( .A(\CARRYB[27][7] ), .B(\ab[28][7] ), .CI(\SUMB[27][8] ), 
        .CO(\CARRYB[28][7] ), .S(\SUMB[28][7] ) );
  FA_X1 S2_27_7 ( .A(\CARRYB[26][7] ), .B(\ab[27][7] ), .CI(\SUMB[26][8] ), 
        .CO(\CARRYB[27][7] ), .S(\SUMB[27][7] ) );
  FA_X1 S2_27_8 ( .A(\CARRYB[26][8] ), .B(\ab[27][8] ), .CI(\SUMB[26][9] ), 
        .CO(\CARRYB[27][8] ), .S(\SUMB[27][8] ) );
  FA_X1 S2_26_8 ( .A(\CARRYB[25][8] ), .B(\ab[26][8] ), .CI(\SUMB[25][9] ), 
        .CO(\CARRYB[26][8] ), .S(\SUMB[26][8] ) );
  FA_X1 S2_26_9 ( .A(\CARRYB[25][9] ), .B(\ab[26][9] ), .CI(\SUMB[25][10] ), 
        .CO(\CARRYB[26][9] ), .S(\SUMB[26][9] ) );
  FA_X1 S2_25_9 ( .A(\CARRYB[24][9] ), .B(\ab[25][9] ), .CI(\SUMB[24][10] ), 
        .CO(\CARRYB[25][9] ), .S(\SUMB[25][9] ) );
  FA_X1 S2_25_10 ( .A(\ab[25][10] ), .B(\CARRYB[24][10] ), .CI(\SUMB[24][11] ), 
        .CO(\CARRYB[25][10] ), .S(\SUMB[25][10] ) );
  FA_X1 S2_24_10 ( .A(\CARRYB[23][10] ), .B(\ab[24][10] ), .CI(\SUMB[23][11] ), 
        .CO(\CARRYB[24][10] ), .S(\SUMB[24][10] ) );
  FA_X1 S2_24_11 ( .A(\CARRYB[23][11] ), .B(\ab[24][11] ), .CI(\SUMB[23][12] ), 
        .CO(\CARRYB[24][11] ), .S(\SUMB[24][11] ) );
  FA_X1 S2_23_11 ( .A(\CARRYB[22][11] ), .B(\ab[23][11] ), .CI(\SUMB[22][12] ), 
        .CO(\CARRYB[23][11] ), .S(\SUMB[23][11] ) );
  FA_X1 S2_23_12 ( .A(\ab[23][12] ), .B(\CARRYB[22][12] ), .CI(\SUMB[22][13] ), 
        .CO(\CARRYB[23][12] ), .S(\SUMB[23][12] ) );
  FA_X1 S2_22_12 ( .A(\CARRYB[21][12] ), .B(\ab[22][12] ), .CI(\SUMB[21][13] ), 
        .CO(\CARRYB[22][12] ), .S(\SUMB[22][12] ) );
  FA_X1 S2_22_13 ( .A(\ab[22][13] ), .B(\CARRYB[21][13] ), .CI(\SUMB[21][14] ), 
        .CO(\CARRYB[22][13] ), .S(\SUMB[22][13] ) );
  FA_X1 S2_21_13 ( .A(\CARRYB[20][13] ), .B(\ab[21][13] ), .CI(\SUMB[20][14] ), 
        .CO(\CARRYB[21][13] ), .S(\SUMB[21][13] ) );
  FA_X1 S2_21_14 ( .A(\ab[21][14] ), .B(\CARRYB[20][14] ), .CI(\SUMB[20][15] ), 
        .CO(\CARRYB[21][14] ), .S(\SUMB[21][14] ) );
  FA_X1 S2_5_29 ( .A(\ab[5][29] ), .B(\CARRYB[4][29] ), .CI(\SUMB[4][30] ), 
        .CO(\CARRYB[5][29] ), .S(\SUMB[5][29] ) );
  FA_X1 S2_7_28 ( .A(\ab[7][28] ), .B(\CARRYB[6][28] ), .CI(\SUMB[6][29] ), 
        .CO(\CARRYB[7][28] ), .S(\SUMB[7][28] ) );
  FA_X1 S2_8_27 ( .A(\ab[8][27] ), .B(\CARRYB[7][27] ), .CI(\SUMB[7][28] ), 
        .CO(\CARRYB[8][27] ), .S(\SUMB[8][27] ) );
  FA_X1 S2_9_26 ( .A(\ab[9][26] ), .B(\CARRYB[8][26] ), .CI(\SUMB[8][27] ), 
        .CO(\CARRYB[9][26] ), .S(\SUMB[9][26] ) );
  FA_X1 S2_10_25 ( .A(\ab[10][25] ), .B(\CARRYB[9][25] ), .CI(\SUMB[9][26] ), 
        .CO(\CARRYB[10][25] ), .S(\SUMB[10][25] ) );
  FA_X1 S2_11_24 ( .A(\ab[11][24] ), .B(\CARRYB[10][24] ), .CI(\SUMB[10][25] ), 
        .CO(\CARRYB[11][24] ), .S(\SUMB[11][24] ) );
  FA_X1 S2_12_23 ( .A(\ab[12][23] ), .B(\CARRYB[11][23] ), .CI(\SUMB[11][24] ), 
        .CO(\CARRYB[12][23] ), .S(\SUMB[12][23] ) );
  FA_X1 S2_13_22 ( .A(\ab[13][22] ), .B(\CARRYB[12][22] ), .CI(\SUMB[12][23] ), 
        .CO(\CARRYB[13][22] ), .S(\SUMB[13][22] ) );
  FA_X1 S2_14_21 ( .A(\ab[14][21] ), .B(\CARRYB[13][21] ), .CI(\SUMB[13][22] ), 
        .CO(\CARRYB[14][21] ), .S(\SUMB[14][21] ) );
  FA_X1 S2_15_20 ( .A(\ab[15][20] ), .B(\CARRYB[14][20] ), .CI(\SUMB[14][21] ), 
        .CO(\CARRYB[15][20] ), .S(\SUMB[15][20] ) );
  FA_X1 S2_16_19 ( .A(\ab[16][19] ), .B(\CARRYB[15][19] ), .CI(\SUMB[15][20] ), 
        .CO(\CARRYB[16][19] ), .S(\SUMB[16][19] ) );
  FA_X1 S2_17_18 ( .A(\ab[17][18] ), .B(\CARRYB[16][18] ), .CI(\SUMB[16][19] ), 
        .CO(\CARRYB[17][18] ), .S(\SUMB[17][18] ) );
  FA_X1 S2_18_17 ( .A(\ab[18][17] ), .B(\CARRYB[17][17] ), .CI(\SUMB[17][18] ), 
        .CO(\CARRYB[18][17] ), .S(\SUMB[18][17] ) );
  FA_X1 S2_19_16 ( .A(\ab[19][16] ), .B(\CARRYB[18][16] ), .CI(\SUMB[18][17] ), 
        .CO(\CARRYB[19][16] ), .S(\SUMB[19][16] ) );
  FA_X1 S2_20_14 ( .A(\ab[20][14] ), .B(\CARRYB[19][14] ), .CI(\SUMB[19][15] ), 
        .CO(\CARRYB[20][14] ), .S(\SUMB[20][14] ) );
  FA_X1 S2_20_15 ( .A(\ab[20][15] ), .B(\CARRYB[19][15] ), .CI(\SUMB[19][16] ), 
        .CO(\CARRYB[20][15] ), .S(\SUMB[20][15] ) );
  FA_X1 S2_17_15 ( .A(\CARRYB[16][15] ), .B(\ab[17][15] ), .CI(\SUMB[16][16] ), 
        .CO(\CARRYB[17][15] ), .S(\SUMB[17][15] ) );
  FA_X1 S2_16_16 ( .A(\CARRYB[15][16] ), .B(\ab[16][16] ), .CI(\SUMB[15][17] ), 
        .CO(\CARRYB[16][16] ), .S(\SUMB[16][16] ) );
  FA_X1 S2_15_17 ( .A(\CARRYB[14][17] ), .B(\ab[15][17] ), .CI(\SUMB[14][18] ), 
        .CO(\CARRYB[15][17] ), .S(\SUMB[15][17] ) );
  FA_X1 S2_14_18 ( .A(\ab[14][18] ), .B(\CARRYB[13][18] ), .CI(\SUMB[13][19] ), 
        .CO(\CARRYB[14][18] ), .S(\SUMB[14][18] ) );
  FA_X1 S2_13_19 ( .A(\CARRYB[12][19] ), .B(\ab[13][19] ), .CI(\SUMB[12][20] ), 
        .CO(\CARRYB[13][19] ), .S(\SUMB[13][19] ) );
  FA_X1 S2_12_20 ( .A(\ab[12][20] ), .B(\CARRYB[11][20] ), .CI(\SUMB[11][21] ), 
        .CO(\CARRYB[12][20] ), .S(\SUMB[12][20] ) );
  FA_X1 S2_11_21 ( .A(\CARRYB[10][21] ), .B(\ab[11][21] ), .CI(\SUMB[10][22] ), 
        .CO(\CARRYB[11][21] ), .S(\SUMB[11][21] ) );
  FA_X1 S2_10_22 ( .A(\ab[10][22] ), .B(\CARRYB[9][22] ), .CI(\SUMB[9][23] ), 
        .CO(\CARRYB[10][22] ), .S(\SUMB[10][22] ) );
  FA_X1 S2_9_23 ( .A(\CARRYB[8][23] ), .B(\ab[9][23] ), .CI(\SUMB[8][24] ), 
        .CO(\CARRYB[9][23] ), .S(\SUMB[9][23] ) );
  FA_X1 S2_8_24 ( .A(\ab[8][24] ), .B(\CARRYB[7][24] ), .CI(\SUMB[7][25] ), 
        .CO(\CARRYB[8][24] ), .S(\SUMB[8][24] ) );
  FA_X1 S2_7_25 ( .A(\CARRYB[6][25] ), .B(\ab[7][25] ), .CI(\SUMB[6][26] ), 
        .CO(\CARRYB[7][25] ), .S(\SUMB[7][25] ) );
  FA_X1 S2_6_26 ( .A(\ab[6][26] ), .B(\CARRYB[5][26] ), .CI(\SUMB[5][27] ), 
        .CO(\CARRYB[6][26] ), .S(\SUMB[6][26] ) );
  FA_X1 S2_5_27 ( .A(\CARRYB[4][27] ), .B(\ab[5][27] ), .CI(\SUMB[4][28] ), 
        .CO(\CARRYB[5][27] ), .S(\SUMB[5][27] ) );
  FA_X1 S2_4_28 ( .A(\ab[4][28] ), .B(\CARRYB[3][28] ), .CI(\SUMB[3][29] ), 
        .CO(\CARRYB[4][28] ), .S(\SUMB[4][28] ) );
  FA_X1 S2_3_29 ( .A(\CARRYB[2][29] ), .B(\ab[3][29] ), .CI(\SUMB[2][30] ), 
        .CO(\CARRYB[3][29] ), .S(\SUMB[3][29] ) );
  FA_X1 S2_6_28 ( .A(\ab[6][28] ), .B(\CARRYB[5][28] ), .CI(\SUMB[5][29] ), 
        .CO(\CARRYB[6][28] ), .S(\SUMB[6][28] ) );
  FA_X1 S2_5_28 ( .A(\CARRYB[4][28] ), .B(\ab[5][28] ), .CI(\SUMB[4][29] ), 
        .CO(\CARRYB[5][28] ), .S(\SUMB[5][28] ) );
  FA_X1 S2_7_27 ( .A(\CARRYB[6][27] ), .B(\ab[7][27] ), .CI(\SUMB[6][28] ), 
        .CO(\CARRYB[7][27] ), .S(\SUMB[7][27] ) );
  FA_X1 S2_6_27 ( .A(\CARRYB[5][27] ), .B(\ab[6][27] ), .CI(\SUMB[5][28] ), 
        .CO(\CARRYB[6][27] ), .S(\SUMB[6][27] ) );
  FA_X1 S2_8_26 ( .A(\ab[8][26] ), .B(\CARRYB[7][26] ), .CI(\SUMB[7][27] ), 
        .CO(\CARRYB[8][26] ), .S(\SUMB[8][26] ) );
  FA_X1 S2_7_26 ( .A(\CARRYB[6][26] ), .B(\ab[7][26] ), .CI(\SUMB[6][27] ), 
        .CO(\CARRYB[7][26] ), .S(\SUMB[7][26] ) );
  FA_X1 S2_9_25 ( .A(\CARRYB[8][25] ), .B(\ab[9][25] ), .CI(\SUMB[8][26] ), 
        .CO(\CARRYB[9][25] ), .S(\SUMB[9][25] ) );
  FA_X1 S2_8_25 ( .A(\CARRYB[7][25] ), .B(\ab[8][25] ), .CI(\SUMB[7][26] ), 
        .CO(\CARRYB[8][25] ), .S(\SUMB[8][25] ) );
  FA_X1 S2_10_24 ( .A(\ab[10][24] ), .B(\CARRYB[9][24] ), .CI(\SUMB[9][25] ), 
        .CO(\CARRYB[10][24] ), .S(\SUMB[10][24] ) );
  FA_X1 S2_9_24 ( .A(\CARRYB[8][24] ), .B(\ab[9][24] ), .CI(\SUMB[8][25] ), 
        .CO(\CARRYB[9][24] ), .S(\SUMB[9][24] ) );
  FA_X1 S2_11_23 ( .A(\CARRYB[10][23] ), .B(\ab[11][23] ), .CI(\SUMB[10][24] ), 
        .CO(\CARRYB[11][23] ), .S(\SUMB[11][23] ) );
  FA_X1 S2_10_23 ( .A(\CARRYB[9][23] ), .B(\ab[10][23] ), .CI(\SUMB[9][24] ), 
        .CO(\CARRYB[10][23] ), .S(\SUMB[10][23] ) );
  FA_X1 S2_12_22 ( .A(\ab[12][22] ), .B(\CARRYB[11][22] ), .CI(\SUMB[11][23] ), 
        .CO(\CARRYB[12][22] ), .S(\SUMB[12][22] ) );
  FA_X1 S2_11_22 ( .A(\ab[11][22] ), .B(\CARRYB[10][22] ), .CI(\SUMB[10][23] ), 
        .CO(\CARRYB[11][22] ), .S(\SUMB[11][22] ) );
  FA_X1 S2_13_21 ( .A(\CARRYB[12][21] ), .B(\ab[13][21] ), .CI(\SUMB[12][22] ), 
        .CO(\CARRYB[13][21] ), .S(\SUMB[13][21] ) );
  FA_X1 S2_12_21 ( .A(\CARRYB[11][21] ), .B(\ab[12][21] ), .CI(\SUMB[11][22] ), 
        .CO(\CARRYB[12][21] ), .S(\SUMB[12][21] ) );
  FA_X1 S2_14_20 ( .A(\ab[14][20] ), .B(\CARRYB[13][20] ), .CI(\SUMB[13][21] ), 
        .CO(\CARRYB[14][20] ), .S(\SUMB[14][20] ) );
  FA_X1 S2_13_20 ( .A(\ab[13][20] ), .B(\CARRYB[12][20] ), .CI(\SUMB[12][21] ), 
        .CO(\CARRYB[13][20] ), .S(\SUMB[13][20] ) );
  FA_X1 S2_15_19 ( .A(\CARRYB[14][19] ), .B(\ab[15][19] ), .CI(\SUMB[14][20] ), 
        .CO(\CARRYB[15][19] ), .S(\SUMB[15][19] ) );
  FA_X1 S2_14_19 ( .A(\CARRYB[13][19] ), .B(\ab[14][19] ), .CI(\SUMB[13][20] ), 
        .CO(\CARRYB[14][19] ), .S(\SUMB[14][19] ) );
  FA_X1 S2_16_18 ( .A(\ab[16][18] ), .B(\CARRYB[15][18] ), .CI(\SUMB[15][19] ), 
        .CO(\CARRYB[16][18] ), .S(\SUMB[16][18] ) );
  FA_X1 S2_15_18 ( .A(\ab[15][18] ), .B(\CARRYB[14][18] ), .CI(\SUMB[14][19] ), 
        .CO(\CARRYB[15][18] ), .S(\SUMB[15][18] ) );
  FA_X1 S2_17_17 ( .A(\CARRYB[16][17] ), .B(\ab[17][17] ), .CI(\SUMB[16][18] ), 
        .CO(\CARRYB[17][17] ), .S(\SUMB[17][17] ) );
  FA_X1 S2_16_17 ( .A(\CARRYB[15][17] ), .B(\ab[16][17] ), .CI(\SUMB[15][18] ), 
        .CO(\CARRYB[16][17] ), .S(\SUMB[16][17] ) );
  FA_X1 S2_18_16 ( .A(\ab[18][16] ), .B(\CARRYB[17][16] ), .CI(\SUMB[17][17] ), 
        .CO(\CARRYB[18][16] ), .S(\SUMB[18][16] ) );
  FA_X1 S2_17_16 ( .A(\ab[17][16] ), .B(\CARRYB[16][16] ), .CI(\SUMB[16][17] ), 
        .CO(\CARRYB[17][16] ), .S(\SUMB[17][16] ) );
  FA_X1 S2_19_14 ( .A(\CARRYB[18][14] ), .B(\ab[19][14] ), .CI(\SUMB[18][15] ), 
        .CO(\CARRYB[19][14] ), .S(\SUMB[19][14] ) );
  FA_X1 S2_19_15 ( .A(\CARRYB[18][15] ), .B(\ab[19][15] ), .CI(\SUMB[18][16] ), 
        .CO(\CARRYB[19][15] ), .S(\SUMB[19][15] ) );
  FA_X1 S2_18_15 ( .A(\CARRYB[17][15] ), .B(\ab[18][15] ), .CI(\SUMB[17][16] ), 
        .CO(\CARRYB[18][15] ), .S(\SUMB[18][15] ) );
  FA_X1 S3_2_30 ( .A(\ab[2][30] ), .B(\ab[1][31] ), .CI(\CARRYB[1][30] ), .CO(
        \CARRYB[2][30] ), .S(\SUMB[2][30] ) );
  INV_X4 U2 ( .A(A[15]), .ZN(n61) );
  CLKBUF_X3 U3 ( .A(n41), .Z(n98) );
  INV_X2 U4 ( .A(B[4]), .ZN(n10) );
  CLKBUF_X2 U5 ( .A(n10), .Z(n176) );
  INV_X2 U6 ( .A(B[2]), .ZN(n14) );
  CLKBUF_X2 U7 ( .A(n14), .Z(n172) );
  INV_X2 U8 ( .A(A[20]), .ZN(n55) );
  INV_X4 U9 ( .A(A[13]), .ZN(n63) );
  INV_X2 U10 ( .A(A[24]), .ZN(n51) );
  INV_X2 U11 ( .A(A[23]), .ZN(n52) );
  INV_X2 U12 ( .A(A[22]), .ZN(n53) );
  INV_X2 U13 ( .A(A[18]), .ZN(n58) );
  INV_X2 U14 ( .A(B[25]), .ZN(n72) );
  CLKBUF_X3 U15 ( .A(n72), .Z(n162) );
  INV_X2 U16 ( .A(A[25]), .ZN(n50) );
  INV_X2 U17 ( .A(A[29]), .ZN(n46) );
  INV_X2 U18 ( .A(A[31]), .ZN(n43) );
  INV_X4 U19 ( .A(A[14]), .ZN(n62) );
  INV_X2 U20 ( .A(A[30]), .ZN(n44) );
  INV_X4 U21 ( .A(A[16]), .ZN(n60) );
  INV_X2 U22 ( .A(A[19]), .ZN(n57) );
  INV_X2 U23 ( .A(A[21]), .ZN(n54) );
  INV_X2 U24 ( .A(A[11]), .ZN(n65) );
  CLKBUF_X3 U25 ( .A(n65), .Z(n92) );
  INV_X2 U26 ( .A(A[28]), .ZN(n47) );
  INV_X2 U27 ( .A(A[27]), .ZN(n48) );
  INV_X2 U28 ( .A(A[12]), .ZN(n64) );
  CLKBUF_X3 U29 ( .A(n64), .Z(n93) );
  INV_X2 U30 ( .A(A[26]), .ZN(n49) );
  INV_X2 U31 ( .A(A[17]), .ZN(n59) );
  CLKBUF_X3 U32 ( .A(n24), .Z(n147) );
  BUF_X2 U33 ( .A(A[0]), .Z(n74) );
  BUF_X1 U34 ( .A(n21), .Z(n156) );
  CLKBUF_X3 U35 ( .A(n67), .Z(net145039) );
  BUF_X2 U36 ( .A(n20), .Z(n159) );
  CLKBUF_X3 U37 ( .A(n15), .Z(n170) );
  INV_X1 U38 ( .A(B[29]), .ZN(n15) );
  INV_X1 U39 ( .A(n81), .ZN(n79) );
  CLKBUF_X3 U40 ( .A(n19), .Z(n161) );
  CLKBUF_X3 U41 ( .A(n23), .Z(n151) );
  XNOR2_X1 U42 ( .A(n73), .B(\ab[0][25] ), .ZN(\SUMB[1][24] ) );
  OR2_X1 U43 ( .A1(n159), .A2(n79), .ZN(n73) );
  AND2_X1 U44 ( .A1(B[27]), .A2(n74), .ZN(\ab[0][27] ) );
  AND2_X1 U45 ( .A1(B[26]), .A2(n74), .ZN(\ab[0][26] ) );
  CLKBUF_X3 U46 ( .A(n27), .Z(n138) );
  INV_X1 U47 ( .A(A[2]), .ZN(n76) );
  INV_X1 U48 ( .A(A[2]), .ZN(n75) );
  CLKBUF_X3 U49 ( .A(n78), .Z(net144717) );
  AND2_X1 U50 ( .A1(B[28]), .A2(n74), .ZN(\ab[0][28] ) );
  CLKBUF_X3 U51 ( .A(net169718), .Z(net144973) );
  CLKBUF_X3 U52 ( .A(n23), .Z(n150) );
  CLKBUF_X2 U53 ( .A(n12), .Z(net144707) );
  CLKBUF_X1 U54 ( .A(B[30]), .Z(n77) );
  CLKBUF_X3 U55 ( .A(n21), .Z(n155) );
  BUF_X1 U56 ( .A(A[1]), .Z(n81) );
  CLKBUF_X3 U57 ( .A(n21), .Z(n157) );
  INV_X1 U58 ( .A(B[30]), .ZN(n78) );
  CLKBUF_X3 U59 ( .A(n67), .Z(net145041) );
  XNOR2_X1 U60 ( .A(\CARRYB[3][29] ), .B(n80), .ZN(\SUMB[4][29] ) );
  XNOR2_X1 U61 ( .A(\SUMB[3][30] ), .B(\ab[4][29] ), .ZN(n80) );
  NAND2_X1 U62 ( .A1(n74), .A2(B[31]), .ZN(net169569) );
  XNOR2_X1 U63 ( .A(n82), .B(\ab[0][26] ), .ZN(\SUMB[1][25] ) );
  OR2_X1 U64 ( .A1(n72), .A2(n56), .ZN(n82) );
  NOR2_X1 U65 ( .A1(n13), .A2(net145037), .ZN(n83) );
  INV_X1 U66 ( .A(n74), .ZN(n84) );
  BUF_X1 U68 ( .A(n67), .Z(net145037) );
  CLKBUF_X1 U70 ( .A(n13), .Z(net144713) );
  AND2_X1 U72 ( .A1(B[28]), .A2(n81), .ZN(\ab[1][28] ) );
  XNOR2_X1 U75 ( .A(n85), .B(n83), .ZN(\SUMB[1][29] ) );
  OR2_X1 U77 ( .A1(n15), .A2(net169718), .ZN(n85) );
  AND2_X1 U79 ( .A1(B[31]), .A2(n81), .ZN(\ab[1][31] ) );
  AND2_X1 U81 ( .A1(B[26]), .A2(n81), .ZN(\ab[1][26] ) );
  AND2_X1 U83 ( .A1(B[28]), .A2(A[2]), .ZN(\ab[2][28] ) );
  NAND2_X1 U85 ( .A1(B[27]), .A2(n81), .ZN(n87) );
  AND2_X1 U87 ( .A1(B[27]), .A2(A[2]), .ZN(\ab[2][27] ) );
  BUF_X1 U89 ( .A(n17), .Z(n165) );
  AND2_X2 U91 ( .A1(\SUMB[31][2] ), .A2(\CARRYB[31][1] ), .ZN(\A2[32] ) );
  AND2_X1 U93 ( .A1(A[2]), .A2(n77), .ZN(\ab[2][30] ) );
  NOR2_X1 U95 ( .A1(n78), .A2(n84), .ZN(\ab[0][30] ) );
  AND2_X1 U97 ( .A1(\ab[1][30] ), .A2(net169256), .ZN(\CARRYB[1][30] ) );
  NOR2_X1 U99 ( .A1(n12), .A2(net145037), .ZN(net169256) );
  INV_X1 U101 ( .A(A[0]), .ZN(n67) );
  INV_X1 U103 ( .A(B[31]), .ZN(n12) );
  CLKBUF_X1 U105 ( .A(n12), .Z(net144709) );
  NOR2_X1 U107 ( .A1(net169827), .A2(net169718), .ZN(\ab[1][30] ) );
  XNOR2_X1 U109 ( .A(\ab[1][30] ), .B(net169569), .ZN(\SUMB[1][30] ) );
  INV_X1 U111 ( .A(A[1]), .ZN(net169718) );
  INV_X1 U113 ( .A(B[30]), .ZN(net169827) );
  INV_X1 U115 ( .A(A[1]), .ZN(n56) );
  INV_X1 U117 ( .A(B[30]), .ZN(n13) );
  NAND2_X1 U119 ( .A1(\CARRYB[3][29] ), .A2(\SUMB[3][30] ), .ZN(net169775) );
  NAND2_X1 U121 ( .A1(\CARRYB[3][29] ), .A2(\ab[4][29] ), .ZN(net169776) );
  NAND2_X1 U123 ( .A1(\CARRYB[2][30] ), .A2(\ab[2][31] ), .ZN(net169226) );
  XNOR2_X1 U125 ( .A(\CARRYB[2][30] ), .B(net169833), .ZN(\SUMB[3][30] ) );
  NAND2_X1 U127 ( .A1(\CARRYB[2][30] ), .A2(\ab[3][30] ), .ZN(net169225) );
  INV_X1 U129 ( .A(A[2]), .ZN(n45) );
  CLKBUF_X2 U131 ( .A(n76), .Z(net144909) );
  CLKBUF_X3 U133 ( .A(net144713), .Z(net169601) );
  AND2_X1 U135 ( .A1(\SUMB[31][4] ), .A2(\CARRYB[31][3] ), .ZN(\A2[34] ) );
  AND2_X1 U137 ( .A1(\SUMB[31][3] ), .A2(\CARRYB[31][2] ), .ZN(\A2[33] ) );
  CLKBUF_X1 U139 ( .A(n17), .Z(n166) );
  CLKBUF_X3 U141 ( .A(n22), .Z(n153) );
  CLKBUF_X1 U143 ( .A(n20), .Z(n160) );
  CLKBUF_X3 U145 ( .A(n20), .Z(n158) );
  XNOR2_X1 U147 ( .A(\ab[3][30] ), .B(\ab[2][31] ), .ZN(net169833) );
  BUF_X1 U149 ( .A(n42), .Z(n94) );
  NAND2_X1 U151 ( .A1(\SUMB[3][30] ), .A2(\ab[4][29] ), .ZN(n86) );
  NAND3_X1 U153 ( .A1(net169775), .A2(net169776), .A3(n86), .ZN(
        \CARRYB[4][29] ) );
  CLKBUF_X1 U155 ( .A(n18), .Z(n164) );
  CLKBUF_X3 U157 ( .A(n18), .Z(n163) );
  CLKBUF_X1 U159 ( .A(n16), .Z(n168) );
  CLKBUF_X3 U161 ( .A(n42), .Z(n95) );
  CLKBUF_X3 U163 ( .A(n42), .Z(n96) );
  XNOR2_X1 U165 ( .A(\ab[0][28] ), .B(n87), .ZN(\SUMB[1][27] ) );
  CLKBUF_X3 U166 ( .A(n17), .Z(n167) );
  CLKBUF_X3 U167 ( .A(n16), .Z(n169) );
  NAND2_X1 U169 ( .A1(\ab[3][30] ), .A2(\ab[2][31] ), .ZN(n88) );
  NAND3_X1 U170 ( .A1(net169225), .A2(net169226), .A3(n88), .ZN(
        \CARRYB[3][30] ) );
  CLKBUF_X1 U171 ( .A(n66), .Z(n91) );
  BUF_X1 U173 ( .A(n26), .Z(n141) );
  BUF_X1 U175 ( .A(n28), .Z(n135) );
  BUF_X1 U177 ( .A(n34), .Z(n117) );
  BUF_X1 U178 ( .A(n29), .Z(n132) );
  BUF_X1 U179 ( .A(n33), .Z(n120) );
  BUF_X1 U181 ( .A(n30), .Z(n129) );
  BUF_X1 U183 ( .A(n32), .Z(n123) );
  BUF_X1 U186 ( .A(n31), .Z(n126) );
  BUF_X1 U188 ( .A(n24), .Z(n146) );
  BUF_X1 U189 ( .A(n26), .Z(n140) );
  BUF_X1 U190 ( .A(n27), .Z(n137) );
  BUF_X1 U191 ( .A(n28), .Z(n134) );
  BUF_X1 U192 ( .A(n29), .Z(n131) );
  BUF_X1 U193 ( .A(n32), .Z(n122) );
  BUF_X1 U194 ( .A(n41), .Z(n97) );
  BUF_X2 U195 ( .A(n22), .Z(n152) );
  BUF_X1 U196 ( .A(n9), .Z(n179) );
  BUF_X1 U197 ( .A(n8), .Z(n182) );
  BUF_X1 U198 ( .A(n7), .Z(n185) );
  BUF_X1 U199 ( .A(n6), .Z(n188) );
  BUF_X1 U200 ( .A(n5), .Z(n191) );
  BUF_X1 U201 ( .A(n35), .Z(n114) );
  BUF_X1 U202 ( .A(n11), .Z(n174) );
  BUF_X1 U203 ( .A(n25), .Z(n144) );
  BUF_X1 U204 ( .A(n4), .Z(n194) );
  BUF_X1 U205 ( .A(n4), .Z(n193) );
  BUF_X1 U206 ( .A(n9), .Z(n178) );
  BUF_X1 U207 ( .A(n30), .Z(n128) );
  BUF_X1 U208 ( .A(n11), .Z(n173) );
  BUF_X1 U209 ( .A(n6), .Z(n187) );
  BUF_X1 U210 ( .A(n5), .Z(n190) );
  BUF_X1 U211 ( .A(n8), .Z(n181) );
  BUF_X1 U212 ( .A(n31), .Z(n125) );
  BUF_X1 U213 ( .A(n7), .Z(n184) );
  BUF_X1 U214 ( .A(n33), .Z(n119) );
  BUF_X1 U215 ( .A(n14), .Z(n171) );
  BUF_X1 U216 ( .A(n35), .Z(n113) );
  BUF_X1 U217 ( .A(n34), .Z(n116) );
  BUF_X1 U218 ( .A(n36), .Z(n111) );
  BUF_X1 U219 ( .A(n25), .Z(n143) );
  BUF_X1 U220 ( .A(n40), .Z(n100) );
  BUF_X1 U221 ( .A(n40), .Z(n99) );
  BUF_X1 U222 ( .A(n39), .Z(n103) );
  BUF_X1 U223 ( .A(n39), .Z(n102) );
  BUF_X1 U224 ( .A(n38), .Z(n106) );
  BUF_X1 U225 ( .A(n38), .Z(n105) );
  BUF_X1 U226 ( .A(n37), .Z(n109) );
  BUF_X1 U227 ( .A(n37), .Z(n108) );
  AND2_X1 U228 ( .A1(\SUMB[31][31] ), .A2(\CARRYB[31][30] ), .ZN(\A2[61] ) );
  AND2_X1 U229 ( .A1(\SUMB[31][7] ), .A2(\CARRYB[31][6] ), .ZN(\A2[37] ) );
  AND2_X1 U230 ( .A1(\SUMB[31][11] ), .A2(\CARRYB[31][10] ), .ZN(\A2[41] ) );
  AND2_X1 U231 ( .A1(\SUMB[31][10] ), .A2(\CARRYB[31][9] ), .ZN(\A2[40] ) );
  AND2_X1 U232 ( .A1(\SUMB[31][5] ), .A2(\CARRYB[31][4] ), .ZN(\A2[35] ) );
  AND2_X1 U233 ( .A1(\SUMB[31][6] ), .A2(\CARRYB[31][5] ), .ZN(\A2[36] ) );
  AND2_X1 U234 ( .A1(\SUMB[31][9] ), .A2(\CARRYB[31][8] ), .ZN(\A2[39] ) );
  AND2_X1 U235 ( .A1(\SUMB[31][13] ), .A2(\CARRYB[31][12] ), .ZN(\A2[43] ) );
  AND2_X1 U236 ( .A1(\SUMB[31][8] ), .A2(\CARRYB[31][7] ), .ZN(\A2[38] ) );
  AND2_X1 U237 ( .A1(\SUMB[31][12] ), .A2(\CARRYB[31][11] ), .ZN(\A2[42] ) );
  AND2_X1 U238 ( .A1(\SUMB[31][14] ), .A2(\CARRYB[31][13] ), .ZN(\A2[44] ) );
  AND2_X1 U239 ( .A1(\SUMB[31][1] ), .A2(\CARRYB[31][0] ), .ZN(\A2[31] ) );
  AND2_X1 U240 ( .A1(\SUMB[31][30] ), .A2(\CARRYB[31][29] ), .ZN(\A2[60] ) );
  AND2_X1 U241 ( .A1(\SUMB[31][24] ), .A2(\CARRYB[31][23] ), .ZN(\A2[54] ) );
  AND2_X1 U242 ( .A1(\SUMB[31][26] ), .A2(\CARRYB[31][25] ), .ZN(\A2[56] ) );
  AND2_X1 U243 ( .A1(\SUMB[31][22] ), .A2(\CARRYB[31][21] ), .ZN(\A2[52] ) );
  AND2_X1 U244 ( .A1(\SUMB[31][20] ), .A2(\CARRYB[31][19] ), .ZN(\A2[50] ) );
  AND2_X1 U245 ( .A1(\SUMB[31][28] ), .A2(\CARRYB[31][27] ), .ZN(\A2[58] ) );
  AND2_X1 U246 ( .A1(\SUMB[31][18] ), .A2(\CARRYB[31][17] ), .ZN(\A2[48] ) );
  AND2_X1 U247 ( .A1(\SUMB[31][15] ), .A2(\CARRYB[31][14] ), .ZN(\A2[45] ) );
  AND2_X1 U248 ( .A1(\SUMB[31][17] ), .A2(\CARRYB[31][16] ), .ZN(\A2[47] ) );
  AND2_X1 U249 ( .A1(\SUMB[31][29] ), .A2(\CARRYB[31][28] ), .ZN(\A2[59] ) );
  AND2_X1 U250 ( .A1(\SUMB[31][25] ), .A2(\CARRYB[31][24] ), .ZN(\A2[55] ) );
  AND2_X1 U251 ( .A1(\SUMB[31][23] ), .A2(\CARRYB[31][22] ), .ZN(\A2[53] ) );
  AND2_X1 U252 ( .A1(\SUMB[31][27] ), .A2(\CARRYB[31][26] ), .ZN(\A2[57] ) );
  AND2_X1 U253 ( .A1(\SUMB[31][21] ), .A2(\CARRYB[31][20] ), .ZN(\A2[51] ) );
  AND2_X1 U254 ( .A1(\SUMB[31][19] ), .A2(\CARRYB[31][18] ), .ZN(\A2[49] ) );
  AND2_X1 U255 ( .A1(\SUMB[31][16] ), .A2(\CARRYB[31][15] ), .ZN(\A2[46] ) );
  NOR2_X1 U256 ( .A1(n15), .A2(n84), .ZN(\ab[0][29] ) );
  NOR2_X1 U257 ( .A1(n72), .A2(net145041), .ZN(\ab[0][25] ) );
  NOR2_X1 U258 ( .A1(n159), .A2(net145039), .ZN(\ab[0][24] ) );
  NOR2_X1 U259 ( .A1(n156), .A2(net145041), .ZN(\ab[0][23] ) );
  NOR2_X1 U260 ( .A1(n151), .A2(net145041), .ZN(\ab[0][21] ) );
  NOR2_X1 U261 ( .A1(n154), .A2(net145039), .ZN(\ab[0][22] ) );
  NOR2_X1 U262 ( .A1(n148), .A2(net145041), .ZN(\ab[0][20] ) );
  NOR2_X1 U263 ( .A1(n142), .A2(net145041), .ZN(\ab[0][19] ) );
  NOR2_X1 U264 ( .A1(n139), .A2(net145039), .ZN(\ab[0][18] ) );
  NOR2_X1 U265 ( .A1(n136), .A2(net145039), .ZN(\ab[0][17] ) );
  NOR2_X1 U266 ( .A1(n133), .A2(net145041), .ZN(\ab[0][16] ) );
  NOR2_X1 U267 ( .A1(n130), .A2(net145039), .ZN(\ab[0][15] ) );
  NOR2_X1 U268 ( .A1(n124), .A2(net145041), .ZN(\ab[0][13] ) );
  NOR2_X1 U269 ( .A1(n127), .A2(net145039), .ZN(\ab[0][14] ) );
  NOR2_X1 U270 ( .A1(n121), .A2(net145039), .ZN(\ab[0][12] ) );
  NOR2_X1 U271 ( .A1(n118), .A2(net145041), .ZN(\ab[0][11] ) );
  NOR2_X1 U272 ( .A1(n115), .A2(net145041), .ZN(\ab[0][10] ) );
  NOR2_X1 U273 ( .A1(n192), .A2(net145039), .ZN(\ab[0][9] ) );
  NOR2_X1 U274 ( .A1(n189), .A2(net145041), .ZN(\ab[0][8] ) );
  NOR2_X1 U275 ( .A1(n186), .A2(net145039), .ZN(\ab[0][7] ) );
  NOR2_X1 U276 ( .A1(n183), .A2(net145039), .ZN(\ab[0][6] ) );
  NOR2_X1 U277 ( .A1(n180), .A2(net145041), .ZN(\ab[0][5] ) );
  NOR2_X1 U278 ( .A1(n177), .A2(net145039), .ZN(\ab[0][4] ) );
  NOR2_X1 U279 ( .A1(n175), .A2(net145041), .ZN(\ab[0][3] ) );
  NOR2_X1 U280 ( .A1(n132), .A2(net144973), .ZN(\ab[1][16] ) );
  NOR2_X1 U281 ( .A1(n129), .A2(net144973), .ZN(\ab[1][15] ) );
  NOR2_X1 U282 ( .A1(n126), .A2(n79), .ZN(\ab[1][14] ) );
  NOR2_X1 U283 ( .A1(n123), .A2(net144973), .ZN(\ab[1][13] ) );
  NOR2_X1 U284 ( .A1(n120), .A2(n79), .ZN(\ab[1][12] ) );
  NOR2_X1 U285 ( .A1(n117), .A2(net144973), .ZN(\ab[1][11] ) );
  NOR2_X1 U286 ( .A1(n114), .A2(n79), .ZN(\ab[1][10] ) );
  NOR2_X1 U287 ( .A1(n173), .A2(n43), .ZN(\ab[31][3] ) );
  NOR2_X1 U288 ( .A1(n176), .A2(n43), .ZN(\ab[31][4] ) );
  NOR2_X1 U289 ( .A1(n184), .A2(n43), .ZN(\ab[31][7] ) );
  NOR2_X1 U290 ( .A1(n187), .A2(n43), .ZN(\ab[31][8] ) );
  NOR2_X1 U291 ( .A1(n116), .A2(n43), .ZN(\ab[31][11] ) );
  NOR2_X1 U292 ( .A1(n119), .A2(n43), .ZN(\ab[31][12] ) );
  NOR2_X1 U293 ( .A1(n178), .A2(n43), .ZN(\ab[31][5] ) );
  NOR2_X1 U294 ( .A1(n181), .A2(n43), .ZN(\ab[31][6] ) );
  NOR2_X1 U295 ( .A1(n113), .A2(n43), .ZN(\ab[31][10] ) );
  NOR2_X1 U296 ( .A1(n190), .A2(n43), .ZN(\ab[31][9] ) );
  NOR2_X1 U297 ( .A1(n122), .A2(n43), .ZN(\ab[31][13] ) );
  NOR2_X1 U298 ( .A1(n125), .A2(n43), .ZN(\ab[31][14] ) );
  NOR2_X1 U299 ( .A1(n128), .A2(n43), .ZN(\ab[31][15] ) );
  NOR2_X1 U300 ( .A1(n131), .A2(n43), .ZN(\ab[31][16] ) );
  NOR2_X1 U301 ( .A1(n165), .A2(n56), .ZN(\ab[1][27] ) );
  NOR2_X1 U302 ( .A1(n161), .A2(net144973), .ZN(\ab[1][25] ) );
  NOR2_X1 U303 ( .A1(n159), .A2(net144973), .ZN(\ab[1][24] ) );
  NOR2_X1 U304 ( .A1(n156), .A2(net144973), .ZN(\ab[1][23] ) );
  NOR2_X1 U305 ( .A1(n153), .A2(net144973), .ZN(\ab[1][22] ) );
  NOR2_X1 U306 ( .A1(n150), .A2(net144973), .ZN(\ab[1][21] ) );
  NOR2_X1 U307 ( .A1(n147), .A2(n79), .ZN(\ab[1][20] ) );
  NOR2_X1 U308 ( .A1(n141), .A2(n56), .ZN(\ab[1][19] ) );
  NOR2_X1 U309 ( .A1(n138), .A2(net144973), .ZN(\ab[1][18] ) );
  NOR2_X1 U310 ( .A1(n135), .A2(net144973), .ZN(\ab[1][17] ) );
  NOR2_X1 U311 ( .A1(n171), .A2(n43), .ZN(\ab[31][2] ) );
  NOR2_X1 U312 ( .A1(n143), .A2(n43), .ZN(\ab[31][1] ) );
  NOR2_X1 U313 ( .A1(n111), .A2(n43), .ZN(\ab[31][0] ) );
  NOR2_X1 U314 ( .A1(n193), .A2(net144709), .ZN(\ab[9][31] ) );
  NOR2_X1 U315 ( .A1(net169601), .A2(n89), .ZN(\ab[10][30] ) );
  NOR2_X1 U316 ( .A1(net144717), .A2(n94), .ZN(\ab[3][30] ) );
  NOR2_X1 U317 ( .A1(net144707), .A2(n45), .ZN(\ab[2][31] ) );
  NOR2_X1 U318 ( .A1(net144709), .A2(n95), .ZN(\ab[3][31] ) );
  NOR2_X1 U319 ( .A1(net144713), .A2(n97), .ZN(\ab[4][30] ) );
  NOR2_X1 U320 ( .A1(net144707), .A2(n97), .ZN(\ab[4][31] ) );
  NOR2_X1 U321 ( .A1(net144717), .A2(n99), .ZN(\ab[5][30] ) );
  NOR2_X1 U322 ( .A1(net144709), .A2(n99), .ZN(\ab[5][31] ) );
  NOR2_X1 U323 ( .A1(net169601), .A2(n102), .ZN(\ab[6][30] ) );
  NOR2_X1 U324 ( .A1(net144707), .A2(n102), .ZN(\ab[6][31] ) );
  NOR2_X1 U325 ( .A1(net144717), .A2(n105), .ZN(\ab[7][30] ) );
  NOR2_X1 U326 ( .A1(net144709), .A2(n105), .ZN(\ab[7][31] ) );
  NOR2_X1 U327 ( .A1(net169601), .A2(n108), .ZN(\ab[8][30] ) );
  NOR2_X1 U328 ( .A1(n193), .A2(net144717), .ZN(\ab[9][30] ) );
  NOR2_X1 U329 ( .A1(net144707), .A2(n108), .ZN(\ab[8][31] ) );
  NOR2_X1 U330 ( .A1(net144707), .A2(n89), .ZN(\ab[10][31] ) );
  NOR2_X1 U331 ( .A1(net169601), .A2(n65), .ZN(\ab[11][30] ) );
  NOR2_X1 U332 ( .A1(net144709), .A2(n65), .ZN(\ab[11][31] ) );
  NOR2_X1 U333 ( .A1(net169601), .A2(n93), .ZN(\ab[12][30] ) );
  NOR2_X1 U334 ( .A1(net144707), .A2(n93), .ZN(\ab[12][31] ) );
  NOR2_X1 U335 ( .A1(net144717), .A2(n63), .ZN(\ab[13][30] ) );
  NOR2_X1 U336 ( .A1(net144717), .A2(n62), .ZN(\ab[14][30] ) );
  NOR2_X1 U337 ( .A1(net144709), .A2(n63), .ZN(\ab[13][31] ) );
  NOR2_X1 U338 ( .A1(net144707), .A2(n62), .ZN(\ab[14][31] ) );
  NOR2_X1 U339 ( .A1(net144717), .A2(n61), .ZN(\ab[15][30] ) );
  NOR2_X1 U340 ( .A1(net144709), .A2(n61), .ZN(\ab[15][31] ) );
  NOR2_X1 U341 ( .A1(net169601), .A2(n60), .ZN(\ab[16][30] ) );
  NOR2_X1 U342 ( .A1(net144707), .A2(n60), .ZN(\ab[16][31] ) );
  NOR2_X1 U343 ( .A1(net144717), .A2(n59), .ZN(\ab[17][30] ) );
  NOR2_X1 U344 ( .A1(n18), .A2(n75), .ZN(\ab[2][26] ) );
  AND2_X1 U345 ( .A1(\ab[1][26] ), .A2(\ab[0][27] ), .ZN(\CARRYB[1][26] ) );
  NOR2_X1 U346 ( .A1(n72), .A2(net144909), .ZN(\ab[2][25] ) );
  AND2_X1 U347 ( .A1(\ab[1][25] ), .A2(\ab[0][26] ), .ZN(\CARRYB[1][25] ) );
  NOR2_X1 U348 ( .A1(n159), .A2(n45), .ZN(\ab[2][24] ) );
  AND2_X1 U349 ( .A1(\ab[1][24] ), .A2(\ab[0][25] ), .ZN(\CARRYB[1][24] ) );
  NOR2_X1 U350 ( .A1(n155), .A2(net144909), .ZN(\ab[2][23] ) );
  AND2_X1 U351 ( .A1(\ab[1][23] ), .A2(\ab[0][24] ), .ZN(\CARRYB[1][23] ) );
  NOR2_X1 U352 ( .A1(n152), .A2(n45), .ZN(\ab[2][22] ) );
  AND2_X1 U353 ( .A1(\ab[1][22] ), .A2(\ab[0][23] ), .ZN(\CARRYB[1][22] ) );
  NOR2_X1 U354 ( .A1(n146), .A2(n45), .ZN(\ab[2][20] ) );
  AND2_X1 U355 ( .A1(\ab[1][20] ), .A2(\ab[0][21] ), .ZN(\CARRYB[1][20] ) );
  NOR2_X1 U356 ( .A1(n137), .A2(n45), .ZN(\ab[2][18] ) );
  AND2_X1 U357 ( .A1(\ab[1][18] ), .A2(\ab[0][19] ), .ZN(\CARRYB[1][18] ) );
  NOR2_X1 U358 ( .A1(n131), .A2(n45), .ZN(\ab[2][16] ) );
  AND2_X1 U359 ( .A1(\ab[1][16] ), .A2(\ab[0][17] ), .ZN(\CARRYB[1][16] ) );
  NOR2_X1 U360 ( .A1(n125), .A2(n45), .ZN(\ab[2][14] ) );
  AND2_X1 U361 ( .A1(\ab[1][14] ), .A2(\ab[0][15] ), .ZN(\CARRYB[1][14] ) );
  NOR2_X1 U362 ( .A1(n119), .A2(n45), .ZN(\ab[2][12] ) );
  AND2_X1 U363 ( .A1(\ab[1][12] ), .A2(\ab[0][13] ), .ZN(\CARRYB[1][12] ) );
  NOR2_X1 U364 ( .A1(n113), .A2(n45), .ZN(\ab[2][10] ) );
  AND2_X1 U365 ( .A1(\ab[1][10] ), .A2(\ab[0][11] ), .ZN(\CARRYB[1][10] ) );
  AND2_X1 U366 ( .A1(\ab[1][29] ), .A2(\ab[0][30] ), .ZN(\CARRYB[1][29] ) );
  NOR2_X1 U367 ( .A1(n15), .A2(n75), .ZN(\ab[2][29] ) );
  AND2_X1 U368 ( .A1(\ab[1][27] ), .A2(\ab[0][28] ), .ZN(\CARRYB[1][27] ) );
  AND2_X1 U369 ( .A1(\ab[1][28] ), .A2(\ab[0][29] ), .ZN(\CARRYB[1][28] ) );
  NOR2_X1 U370 ( .A1(n187), .A2(n45), .ZN(\ab[2][8] ) );
  AND2_X1 U371 ( .A1(\ab[1][8] ), .A2(\ab[0][9] ), .ZN(\CARRYB[1][8] ) );
  NOR2_X1 U372 ( .A1(n181), .A2(n45), .ZN(\ab[2][6] ) );
  AND2_X1 U373 ( .A1(\ab[1][6] ), .A2(\ab[0][7] ), .ZN(\CARRYB[1][6] ) );
  NOR2_X1 U374 ( .A1(n176), .A2(n45), .ZN(\ab[2][4] ) );
  AND2_X1 U375 ( .A1(\ab[1][4] ), .A2(\ab[0][5] ), .ZN(\CARRYB[1][4] ) );
  NOR2_X1 U376 ( .A1(n176), .A2(n44), .ZN(\ab[30][4] ) );
  NOR2_X1 U377 ( .A1(n187), .A2(n44), .ZN(\ab[30][8] ) );
  NOR2_X1 U378 ( .A1(n184), .A2(n44), .ZN(\ab[30][7] ) );
  NOR2_X1 U379 ( .A1(n190), .A2(n44), .ZN(\ab[30][9] ) );
  NOR2_X1 U380 ( .A1(n119), .A2(n44), .ZN(\ab[30][12] ) );
  NOR2_X1 U381 ( .A1(n181), .A2(n44), .ZN(\ab[30][6] ) );
  NOR2_X1 U382 ( .A1(n113), .A2(n44), .ZN(\ab[30][10] ) );
  NOR2_X1 U383 ( .A1(n122), .A2(n44), .ZN(\ab[30][13] ) );
  NOR2_X1 U384 ( .A1(n176), .A2(n46), .ZN(\ab[29][4] ) );
  NOR2_X1 U385 ( .A1(n178), .A2(n46), .ZN(\ab[29][5] ) );
  NOR2_X1 U386 ( .A1(n187), .A2(n46), .ZN(\ab[29][8] ) );
  NOR2_X1 U387 ( .A1(n181), .A2(n46), .ZN(\ab[29][6] ) );
  NOR2_X1 U388 ( .A1(n125), .A2(n44), .ZN(\ab[30][14] ) );
  NOR2_X1 U389 ( .A1(n184), .A2(n46), .ZN(\ab[29][7] ) );
  NOR2_X1 U390 ( .A1(n113), .A2(n46), .ZN(\ab[29][10] ) );
  NOR2_X1 U391 ( .A1(n119), .A2(n46), .ZN(\ab[29][12] ) );
  NOR2_X1 U392 ( .A1(n116), .A2(n46), .ZN(\ab[29][11] ) );
  NOR2_X1 U393 ( .A1(n128), .A2(n44), .ZN(\ab[30][15] ) );
  NOR2_X1 U394 ( .A1(n122), .A2(n46), .ZN(\ab[29][13] ) );
  NOR2_X1 U395 ( .A1(n178), .A2(n47), .ZN(\ab[28][5] ) );
  NOR2_X1 U396 ( .A1(n131), .A2(n44), .ZN(\ab[30][16] ) );
  NOR2_X1 U397 ( .A1(n176), .A2(n47), .ZN(\ab[28][4] ) );
  NOR2_X1 U398 ( .A1(n181), .A2(n47), .ZN(\ab[28][6] ) );
  NOR2_X1 U399 ( .A1(n190), .A2(n47), .ZN(\ab[28][9] ) );
  NOR2_X1 U400 ( .A1(n125), .A2(n46), .ZN(\ab[29][14] ) );
  NOR2_X1 U401 ( .A1(n187), .A2(n47), .ZN(\ab[28][8] ) );
  NOR2_X1 U402 ( .A1(n184), .A2(n47), .ZN(\ab[28][7] ) );
  NOR2_X1 U403 ( .A1(n113), .A2(n47), .ZN(\ab[28][10] ) );
  NOR2_X1 U404 ( .A1(n134), .A2(n44), .ZN(\ab[30][17] ) );
  NOR2_X1 U405 ( .A1(n167), .A2(n98), .ZN(\ab[4][27] ) );
  NOR2_X1 U406 ( .A1(n166), .A2(n100), .ZN(\ab[5][27] ) );
  NOR2_X1 U407 ( .A1(n162), .A2(n103), .ZN(\ab[6][25] ) );
  NOR2_X1 U408 ( .A1(n161), .A2(n106), .ZN(\ab[7][25] ) );
  NOR2_X1 U409 ( .A1(n72), .A2(n109), .ZN(\ab[8][25] ) );
  NOR2_X1 U410 ( .A1(n155), .A2(n90), .ZN(\ab[10][23] ) );
  NOR2_X1 U411 ( .A1(n150), .A2(n64), .ZN(\ab[12][21] ) );
  NOR2_X1 U412 ( .A1(n142), .A2(n62), .ZN(\ab[14][19] ) );
  NOR2_X1 U413 ( .A1(n185), .A2(n50), .ZN(\ab[25][7] ) );
  NOR2_X1 U414 ( .A1(n136), .A2(n60), .ZN(\ab[16][17] ) );
  NOR2_X1 U415 ( .A1(n129), .A2(n58), .ZN(\ab[18][15] ) );
  NOR2_X1 U416 ( .A1(n123), .A2(n55), .ZN(\ab[20][13] ) );
  NOR2_X1 U417 ( .A1(n117), .A2(n53), .ZN(\ab[22][11] ) );
  NOR2_X1 U418 ( .A1(n191), .A2(n51), .ZN(\ab[24][9] ) );
  NOR2_X1 U419 ( .A1(n185), .A2(n49), .ZN(\ab[26][7] ) );
  NOR2_X1 U420 ( .A1(n170), .A2(n94), .ZN(\ab[3][29] ) );
  NOR2_X1 U421 ( .A1(n167), .A2(n103), .ZN(\ab[6][27] ) );
  NOR2_X1 U422 ( .A1(n170), .A2(n97), .ZN(\ab[4][29] ) );
  NOR2_X1 U423 ( .A1(n155), .A2(n92), .ZN(\ab[11][23] ) );
  NOR2_X1 U424 ( .A1(n151), .A2(n63), .ZN(\ab[13][21] ) );
  NOR2_X1 U425 ( .A1(n142), .A2(n61), .ZN(\ab[15][19] ) );
  NOR2_X1 U426 ( .A1(n135), .A2(n59), .ZN(\ab[17][17] ) );
  NOR2_X1 U427 ( .A1(n129), .A2(n57), .ZN(\ab[19][15] ) );
  NOR2_X1 U428 ( .A1(n123), .A2(n54), .ZN(\ab[21][13] ) );
  NOR2_X1 U429 ( .A1(n117), .A2(n52), .ZN(\ab[23][11] ) );
  NOR2_X1 U430 ( .A1(n191), .A2(n50), .ZN(\ab[25][9] ) );
  NOR2_X1 U431 ( .A1(n185), .A2(n48), .ZN(\ab[27][7] ) );
  NOR2_X1 U432 ( .A1(n194), .A2(n162), .ZN(\ab[9][25] ) );
  NOR2_X1 U433 ( .A1(n166), .A2(n106), .ZN(\ab[7][27] ) );
  NOR2_X1 U434 ( .A1(n170), .A2(n99), .ZN(\ab[5][29] ) );
  NOR2_X1 U435 ( .A1(n149), .A2(n62), .ZN(\ab[14][21] ) );
  NOR2_X1 U436 ( .A1(n142), .A2(n60), .ZN(\ab[16][19] ) );
  NOR2_X1 U437 ( .A1(n135), .A2(n58), .ZN(\ab[18][17] ) );
  NOR2_X1 U438 ( .A1(n129), .A2(n55), .ZN(\ab[20][15] ) );
  NOR2_X1 U439 ( .A1(n123), .A2(n53), .ZN(\ab[22][13] ) );
  NOR2_X1 U440 ( .A1(n117), .A2(n51), .ZN(\ab[24][11] ) );
  NOR2_X1 U441 ( .A1(n191), .A2(n49), .ZN(\ab[26][9] ) );
  NOR2_X1 U442 ( .A1(n155), .A2(n64), .ZN(\ab[12][23] ) );
  NOR2_X1 U443 ( .A1(n161), .A2(n90), .ZN(\ab[10][25] ) );
  NOR2_X1 U444 ( .A1(n167), .A2(n109), .ZN(\ab[8][27] ) );
  NOR2_X1 U445 ( .A1(n170), .A2(n102), .ZN(\ab[6][29] ) );
  NOR2_X1 U446 ( .A1(n164), .A2(n106), .ZN(\ab[7][26] ) );
  NOR2_X1 U447 ( .A1(n194), .A2(n160), .ZN(\ab[9][24] ) );
  NOR2_X1 U448 ( .A1(n154), .A2(n92), .ZN(\ab[11][22] ) );
  NOR2_X1 U449 ( .A1(n148), .A2(n63), .ZN(\ab[13][20] ) );
  NOR2_X1 U450 ( .A1(n139), .A2(n61), .ZN(\ab[15][18] ) );
  NOR2_X1 U451 ( .A1(n132), .A2(n59), .ZN(\ab[17][16] ) );
  NOR2_X1 U452 ( .A1(n126), .A2(n57), .ZN(\ab[19][14] ) );
  NOR2_X1 U453 ( .A1(n120), .A2(n54), .ZN(\ab[21][12] ) );
  NOR2_X1 U454 ( .A1(n114), .A2(n52), .ZN(\ab[23][10] ) );
  NOR2_X1 U455 ( .A1(n188), .A2(n50), .ZN(\ab[25][8] ) );
  NOR2_X1 U456 ( .A1(n182), .A2(n48), .ZN(\ab[27][6] ) );
  NOR2_X1 U457 ( .A1(n169), .A2(n99), .ZN(\ab[5][28] ) );
  NOR2_X1 U458 ( .A1(n158), .A2(n90), .ZN(\ab[10][24] ) );
  NOR2_X1 U459 ( .A1(n154), .A2(n64), .ZN(\ab[12][22] ) );
  NOR2_X1 U460 ( .A1(n148), .A2(n62), .ZN(\ab[14][20] ) );
  NOR2_X1 U461 ( .A1(n139), .A2(n60), .ZN(\ab[16][18] ) );
  NOR2_X1 U462 ( .A1(n132), .A2(n58), .ZN(\ab[18][16] ) );
  NOR2_X1 U463 ( .A1(n126), .A2(n55), .ZN(\ab[20][14] ) );
  NOR2_X1 U464 ( .A1(n120), .A2(n53), .ZN(\ab[22][12] ) );
  NOR2_X1 U465 ( .A1(n114), .A2(n51), .ZN(\ab[24][10] ) );
  NOR2_X1 U466 ( .A1(n163), .A2(n109), .ZN(\ab[8][26] ) );
  NOR2_X1 U467 ( .A1(n188), .A2(n49), .ZN(\ab[26][8] ) );
  NOR2_X1 U468 ( .A1(n168), .A2(n102), .ZN(\ab[6][28] ) );
  NOR2_X1 U469 ( .A1(n154), .A2(n63), .ZN(\ab[13][22] ) );
  NOR2_X1 U470 ( .A1(n148), .A2(n61), .ZN(\ab[15][20] ) );
  NOR2_X1 U471 ( .A1(n138), .A2(n59), .ZN(\ab[17][18] ) );
  NOR2_X1 U472 ( .A1(n132), .A2(n57), .ZN(\ab[19][16] ) );
  NOR2_X1 U473 ( .A1(n126), .A2(n54), .ZN(\ab[21][14] ) );
  NOR2_X1 U474 ( .A1(n120), .A2(n52), .ZN(\ab[23][12] ) );
  NOR2_X1 U475 ( .A1(n114), .A2(n50), .ZN(\ab[25][10] ) );
  NOR2_X1 U476 ( .A1(n188), .A2(n48), .ZN(\ab[27][8] ) );
  NOR2_X1 U477 ( .A1(n148), .A2(n60), .ZN(\ab[16][20] ) );
  NOR2_X1 U478 ( .A1(n138), .A2(n58), .ZN(\ab[18][18] ) );
  NOR2_X1 U479 ( .A1(n132), .A2(n55), .ZN(\ab[20][16] ) );
  NOR2_X1 U480 ( .A1(n126), .A2(n53), .ZN(\ab[22][14] ) );
  NOR2_X1 U481 ( .A1(n120), .A2(n51), .ZN(\ab[24][12] ) );
  NOR2_X1 U482 ( .A1(n114), .A2(n49), .ZN(\ab[26][10] ) );
  NOR2_X1 U483 ( .A1(n160), .A2(n92), .ZN(\ab[11][24] ) );
  NOR2_X1 U484 ( .A1(n154), .A2(n62), .ZN(\ab[14][22] ) );
  NOR2_X1 U485 ( .A1(n194), .A2(n164), .ZN(\ab[9][26] ) );
  NOR2_X1 U486 ( .A1(n158), .A2(n64), .ZN(\ab[12][24] ) );
  NOR2_X1 U487 ( .A1(n169), .A2(n105), .ZN(\ab[7][28] ) );
  NOR2_X1 U488 ( .A1(n163), .A2(n90), .ZN(\ab[10][26] ) );
  NOR2_X1 U489 ( .A1(n168), .A2(n108), .ZN(\ab[8][28] ) );
  NOR2_X1 U490 ( .A1(n169), .A2(n97), .ZN(\ab[4][28] ) );
  NOR2_X1 U491 ( .A1(n164), .A2(n103), .ZN(\ab[6][26] ) );
  NOR2_X1 U492 ( .A1(n158), .A2(n109), .ZN(\ab[8][24] ) );
  NOR2_X1 U493 ( .A1(n154), .A2(n90), .ZN(\ab[10][22] ) );
  NOR2_X1 U494 ( .A1(n148), .A2(n64), .ZN(\ab[12][20] ) );
  NOR2_X1 U495 ( .A1(n139), .A2(n62), .ZN(\ab[14][18] ) );
  NOR2_X1 U496 ( .A1(n133), .A2(n60), .ZN(\ab[16][16] ) );
  NOR2_X1 U497 ( .A1(n126), .A2(n58), .ZN(\ab[18][14] ) );
  NOR2_X1 U498 ( .A1(n120), .A2(n55), .ZN(\ab[20][12] ) );
  NOR2_X1 U499 ( .A1(n114), .A2(n53), .ZN(\ab[22][10] ) );
  NOR2_X1 U500 ( .A1(n188), .A2(n51), .ZN(\ab[24][8] ) );
  NOR2_X1 U501 ( .A1(n182), .A2(n49), .ZN(\ab[26][6] ) );
  NOR2_X1 U502 ( .A1(n168), .A2(n94), .ZN(\ab[3][28] ) );
  NOR2_X1 U503 ( .A1(n163), .A2(n100), .ZN(\ab[5][26] ) );
  NOR2_X1 U504 ( .A1(n160), .A2(n106), .ZN(\ab[7][24] ) );
  NOR2_X1 U505 ( .A1(n194), .A2(n152), .ZN(\ab[9][22] ) );
  NOR2_X1 U506 ( .A1(n148), .A2(n92), .ZN(\ab[11][20] ) );
  NOR2_X1 U507 ( .A1(n139), .A2(n63), .ZN(\ab[13][18] ) );
  NOR2_X1 U508 ( .A1(n133), .A2(n61), .ZN(\ab[15][16] ) );
  NOR2_X1 U509 ( .A1(n126), .A2(n59), .ZN(\ab[17][14] ) );
  NOR2_X1 U510 ( .A1(n120), .A2(n57), .ZN(\ab[19][12] ) );
  NOR2_X1 U511 ( .A1(n114), .A2(n54), .ZN(\ab[21][10] ) );
  NOR2_X1 U512 ( .A1(n188), .A2(n52), .ZN(\ab[23][8] ) );
  NOR2_X1 U513 ( .A1(n182), .A2(n50), .ZN(\ab[25][6] ) );
  NOR2_X1 U514 ( .A1(n10), .A2(n48), .ZN(\ab[27][4] ) );
  NOR2_X1 U515 ( .A1(n141), .A2(n59), .ZN(\ab[17][19] ) );
  NOR2_X1 U516 ( .A1(n135), .A2(n57), .ZN(\ab[19][17] ) );
  NOR2_X1 U517 ( .A1(n129), .A2(n54), .ZN(\ab[21][15] ) );
  NOR2_X1 U518 ( .A1(n123), .A2(n52), .ZN(\ab[23][13] ) );
  NOR2_X1 U519 ( .A1(n117), .A2(n50), .ZN(\ab[25][11] ) );
  NOR2_X1 U520 ( .A1(n191), .A2(n48), .ZN(\ab[27][9] ) );
  NOR2_X1 U521 ( .A1(n150), .A2(n61), .ZN(\ab[15][21] ) );
  NOR2_X1 U522 ( .A1(n157), .A2(n63), .ZN(\ab[13][23] ) );
  NOR2_X1 U523 ( .A1(n72), .A2(n92), .ZN(\ab[11][25] ) );
  NOR2_X1 U524 ( .A1(n194), .A2(n166), .ZN(\ab[9][27] ) );
  NOR2_X1 U525 ( .A1(n170), .A2(n105), .ZN(\ab[7][29] ) );
  NOR2_X1 U526 ( .A1(n116), .A2(n47), .ZN(\ab[28][11] ) );
  NOR2_X1 U527 ( .A1(n161), .A2(n98), .ZN(\ab[4][25] ) );
  NOR2_X1 U528 ( .A1(n72), .A2(n100), .ZN(\ab[5][25] ) );
  NOR2_X1 U529 ( .A1(n157), .A2(n106), .ZN(\ab[7][23] ) );
  NOR2_X1 U530 ( .A1(n166), .A2(n95), .ZN(\ab[3][27] ) );
  NOR2_X1 U531 ( .A1(n163), .A2(n98), .ZN(\ab[4][26] ) );
  NOR2_X1 U532 ( .A1(n160), .A2(n103), .ZN(\ab[6][24] ) );
  NOR2_X1 U533 ( .A1(n152), .A2(n109), .ZN(\ab[8][22] ) );
  NOR2_X1 U534 ( .A1(n148), .A2(n90), .ZN(\ab[10][20] ) );
  NOR2_X1 U535 ( .A1(n139), .A2(n64), .ZN(\ab[12][18] ) );
  NOR2_X1 U536 ( .A1(n133), .A2(n62), .ZN(\ab[14][16] ) );
  NOR2_X1 U537 ( .A1(n127), .A2(n60), .ZN(\ab[16][14] ) );
  NOR2_X1 U538 ( .A1(n120), .A2(n58), .ZN(\ab[18][12] ) );
  NOR2_X1 U539 ( .A1(n114), .A2(n55), .ZN(\ab[20][10] ) );
  NOR2_X1 U540 ( .A1(n188), .A2(n53), .ZN(\ab[22][8] ) );
  NOR2_X1 U541 ( .A1(n182), .A2(n51), .ZN(\ab[24][6] ) );
  NOR2_X1 U542 ( .A1(n10), .A2(n49), .ZN(\ab[26][4] ) );
  NOR2_X1 U543 ( .A1(n158), .A2(n100), .ZN(\ab[5][24] ) );
  NOR2_X1 U544 ( .A1(n152), .A2(n106), .ZN(\ab[7][22] ) );
  NOR2_X1 U545 ( .A1(n194), .A2(n146), .ZN(\ab[9][20] ) );
  NOR2_X1 U546 ( .A1(n139), .A2(n92), .ZN(\ab[11][18] ) );
  NOR2_X1 U547 ( .A1(n133), .A2(n63), .ZN(\ab[13][16] ) );
  NOR2_X1 U548 ( .A1(n127), .A2(n61), .ZN(\ab[15][14] ) );
  NOR2_X1 U549 ( .A1(n120), .A2(n59), .ZN(\ab[17][12] ) );
  NOR2_X1 U550 ( .A1(n164), .A2(n96), .ZN(\ab[3][26] ) );
  NOR2_X1 U551 ( .A1(n114), .A2(n57), .ZN(\ab[19][10] ) );
  NOR2_X1 U552 ( .A1(n188), .A2(n54), .ZN(\ab[21][8] ) );
  NOR2_X1 U553 ( .A1(n182), .A2(n52), .ZN(\ab[23][6] ) );
  NOR2_X1 U554 ( .A1(n10), .A2(n50), .ZN(\ab[25][4] ) );
  NOR2_X1 U555 ( .A1(n135), .A2(n55), .ZN(\ab[20][17] ) );
  NOR2_X1 U556 ( .A1(n129), .A2(n53), .ZN(\ab[22][15] ) );
  NOR2_X1 U557 ( .A1(n123), .A2(n51), .ZN(\ab[24][13] ) );
  NOR2_X1 U558 ( .A1(n117), .A2(n49), .ZN(\ab[26][11] ) );
  NOR2_X1 U559 ( .A1(n141), .A2(n58), .ZN(\ab[18][19] ) );
  NOR2_X1 U560 ( .A1(n151), .A2(n60), .ZN(\ab[16][21] ) );
  NOR2_X1 U561 ( .A1(n157), .A2(n62), .ZN(\ab[14][23] ) );
  NOR2_X1 U562 ( .A1(n162), .A2(n64), .ZN(\ab[12][25] ) );
  NOR2_X1 U563 ( .A1(n167), .A2(n90), .ZN(\ab[10][27] ) );
  NOR2_X1 U564 ( .A1(n170), .A2(n108), .ZN(\ab[8][29] ) );
  NOR2_X1 U565 ( .A1(n158), .A2(n98), .ZN(\ab[4][24] ) );
  NOR2_X1 U566 ( .A1(n152), .A2(n103), .ZN(\ab[6][22] ) );
  NOR2_X1 U567 ( .A1(n146), .A2(n109), .ZN(\ab[8][20] ) );
  NOR2_X1 U568 ( .A1(n139), .A2(n90), .ZN(\ab[10][18] ) );
  NOR2_X1 U569 ( .A1(n133), .A2(n93), .ZN(\ab[12][16] ) );
  NOR2_X1 U570 ( .A1(n127), .A2(n62), .ZN(\ab[14][14] ) );
  NOR2_X1 U571 ( .A1(n121), .A2(n60), .ZN(\ab[16][12] ) );
  NOR2_X1 U572 ( .A1(n114), .A2(n58), .ZN(\ab[18][10] ) );
  NOR2_X1 U573 ( .A1(n188), .A2(n55), .ZN(\ab[20][8] ) );
  NOR2_X1 U574 ( .A1(n182), .A2(n53), .ZN(\ab[22][6] ) );
  NOR2_X1 U575 ( .A1(n10), .A2(n51), .ZN(\ab[24][4] ) );
  NOR2_X1 U576 ( .A1(n147), .A2(n59), .ZN(\ab[17][20] ) );
  NOR2_X1 U577 ( .A1(n138), .A2(n57), .ZN(\ab[19][18] ) );
  NOR2_X1 U578 ( .A1(n132), .A2(n54), .ZN(\ab[21][16] ) );
  NOR2_X1 U579 ( .A1(n126), .A2(n52), .ZN(\ab[23][14] ) );
  NOR2_X1 U580 ( .A1(n120), .A2(n50), .ZN(\ab[25][12] ) );
  NOR2_X1 U581 ( .A1(n154), .A2(n61), .ZN(\ab[15][22] ) );
  NOR2_X1 U582 ( .A1(n114), .A2(n48), .ZN(\ab[27][10] ) );
  NOR2_X1 U583 ( .A1(n158), .A2(n63), .ZN(\ab[13][24] ) );
  NOR2_X1 U584 ( .A1(n164), .A2(n92), .ZN(\ab[11][26] ) );
  NOR2_X1 U585 ( .A1(n193), .A2(n169), .ZN(\ab[9][28] ) );
  NOR2_X1 U586 ( .A1(n129), .A2(n52), .ZN(\ab[23][15] ) );
  NOR2_X1 U587 ( .A1(n123), .A2(n50), .ZN(\ab[25][13] ) );
  NOR2_X1 U588 ( .A1(n117), .A2(n48), .ZN(\ab[27][11] ) );
  NOR2_X1 U589 ( .A1(n135), .A2(n54), .ZN(\ab[21][17] ) );
  NOR2_X1 U590 ( .A1(n141), .A2(n57), .ZN(\ab[19][19] ) );
  NOR2_X1 U591 ( .A1(n149), .A2(n59), .ZN(\ab[17][21] ) );
  NOR2_X1 U592 ( .A1(n157), .A2(n61), .ZN(\ab[15][23] ) );
  NOR2_X1 U593 ( .A1(n161), .A2(n63), .ZN(\ab[13][25] ) );
  NOR2_X1 U594 ( .A1(n167), .A2(n92), .ZN(\ab[11][27] ) );
  NOR2_X1 U595 ( .A1(n193), .A2(n170), .ZN(\ab[9][29] ) );
  NOR2_X1 U596 ( .A1(n160), .A2(n96), .ZN(\ab[3][24] ) );
  NOR2_X1 U597 ( .A1(n152), .A2(n100), .ZN(\ab[5][22] ) );
  NOR2_X1 U598 ( .A1(n146), .A2(n106), .ZN(\ab[7][20] ) );
  NOR2_X1 U599 ( .A1(n194), .A2(n137), .ZN(\ab[9][18] ) );
  NOR2_X1 U600 ( .A1(n133), .A2(n92), .ZN(\ab[11][16] ) );
  NOR2_X1 U601 ( .A1(n127), .A2(n63), .ZN(\ab[13][14] ) );
  NOR2_X1 U602 ( .A1(n121), .A2(n61), .ZN(\ab[15][12] ) );
  NOR2_X1 U603 ( .A1(n114), .A2(n59), .ZN(\ab[17][10] ) );
  NOR2_X1 U604 ( .A1(n188), .A2(n57), .ZN(\ab[19][8] ) );
  NOR2_X1 U605 ( .A1(n182), .A2(n54), .ZN(\ab[21][6] ) );
  NOR2_X1 U606 ( .A1(n10), .A2(n52), .ZN(\ab[23][4] ) );
  NOR2_X1 U607 ( .A1(n128), .A2(n46), .ZN(\ab[29][15] ) );
  NOR2_X1 U608 ( .A1(n132), .A2(n53), .ZN(\ab[22][16] ) );
  NOR2_X1 U609 ( .A1(n126), .A2(n51), .ZN(\ab[24][14] ) );
  NOR2_X1 U610 ( .A1(n120), .A2(n49), .ZN(\ab[26][12] ) );
  NOR2_X1 U611 ( .A1(n138), .A2(n55), .ZN(\ab[20][18] ) );
  NOR2_X1 U612 ( .A1(n147), .A2(n58), .ZN(\ab[18][20] ) );
  NOR2_X1 U613 ( .A1(n154), .A2(n60), .ZN(\ab[16][22] ) );
  NOR2_X1 U614 ( .A1(n160), .A2(n62), .ZN(\ab[14][24] ) );
  NOR2_X1 U615 ( .A1(n163), .A2(n64), .ZN(\ab[12][26] ) );
  NOR2_X1 U616 ( .A1(n168), .A2(n89), .ZN(\ab[10][28] ) );
  NOR2_X1 U617 ( .A1(n119), .A2(n47), .ZN(\ab[28][12] ) );
  NOR2_X1 U618 ( .A1(n126), .A2(n50), .ZN(\ab[25][14] ) );
  NOR2_X1 U619 ( .A1(n120), .A2(n48), .ZN(\ab[27][12] ) );
  NOR2_X1 U620 ( .A1(n132), .A2(n52), .ZN(\ab[23][16] ) );
  NOR2_X1 U621 ( .A1(n138), .A2(n54), .ZN(\ab[21][18] ) );
  NOR2_X1 U622 ( .A1(n147), .A2(n57), .ZN(\ab[19][20] ) );
  NOR2_X1 U623 ( .A1(n153), .A2(n59), .ZN(\ab[17][22] ) );
  NOR2_X1 U624 ( .A1(n158), .A2(n61), .ZN(\ab[15][24] ) );
  NOR2_X1 U625 ( .A1(n163), .A2(n63), .ZN(\ab[13][26] ) );
  NOR2_X1 U626 ( .A1(n168), .A2(n65), .ZN(\ab[11][28] ) );
  NOR2_X1 U627 ( .A1(n149), .A2(n100), .ZN(\ab[5][21] ) );
  NOR2_X1 U628 ( .A1(n123), .A2(n49), .ZN(\ab[26][13] ) );
  NOR2_X1 U629 ( .A1(n129), .A2(n51), .ZN(\ab[24][15] ) );
  NOR2_X1 U630 ( .A1(n135), .A2(n53), .ZN(\ab[22][17] ) );
  NOR2_X1 U631 ( .A1(n141), .A2(n55), .ZN(\ab[20][19] ) );
  NOR2_X1 U632 ( .A1(n150), .A2(n58), .ZN(\ab[18][21] ) );
  NOR2_X1 U633 ( .A1(n155), .A2(n60), .ZN(\ab[16][23] ) );
  NOR2_X1 U634 ( .A1(n72), .A2(n62), .ZN(\ab[14][25] ) );
  NOR2_X1 U635 ( .A1(n167), .A2(n64), .ZN(\ab[12][27] ) );
  NOR2_X1 U636 ( .A1(n170), .A2(n89), .ZN(\ab[10][29] ) );
  NOR2_X1 U637 ( .A1(n152), .A2(n98), .ZN(\ab[4][22] ) );
  NOR2_X1 U638 ( .A1(n146), .A2(n103), .ZN(\ab[6][20] ) );
  NOR2_X1 U639 ( .A1(n137), .A2(n109), .ZN(\ab[8][18] ) );
  NOR2_X1 U640 ( .A1(n133), .A2(n91), .ZN(\ab[10][16] ) );
  NOR2_X1 U641 ( .A1(n127), .A2(n64), .ZN(\ab[12][14] ) );
  NOR2_X1 U642 ( .A1(n121), .A2(n62), .ZN(\ab[14][12] ) );
  NOR2_X1 U643 ( .A1(n115), .A2(n60), .ZN(\ab[16][10] ) );
  NOR2_X1 U644 ( .A1(n188), .A2(n58), .ZN(\ab[18][8] ) );
  NOR2_X1 U645 ( .A1(n182), .A2(n55), .ZN(\ab[20][6] ) );
  NOR2_X1 U646 ( .A1(n10), .A2(n53), .ZN(\ab[22][4] ) );
  NOR2_X1 U647 ( .A1(n152), .A2(n95), .ZN(\ab[3][22] ) );
  NOR2_X1 U648 ( .A1(n146), .A2(n100), .ZN(\ab[5][20] ) );
  NOR2_X1 U649 ( .A1(n137), .A2(n106), .ZN(\ab[7][18] ) );
  NOR2_X1 U650 ( .A1(n195), .A2(n131), .ZN(\ab[9][16] ) );
  NOR2_X1 U651 ( .A1(n127), .A2(n65), .ZN(\ab[11][14] ) );
  NOR2_X1 U652 ( .A1(n121), .A2(n63), .ZN(\ab[13][12] ) );
  NOR2_X1 U653 ( .A1(n115), .A2(n61), .ZN(\ab[15][10] ) );
  NOR2_X1 U654 ( .A1(n188), .A2(n59), .ZN(\ab[17][8] ) );
  NOR2_X1 U655 ( .A1(n182), .A2(n57), .ZN(\ab[19][6] ) );
  NOR2_X1 U656 ( .A1(n10), .A2(n54), .ZN(\ab[21][4] ) );
  NOR2_X1 U657 ( .A1(n122), .A2(n47), .ZN(\ab[28][13] ) );
  NOR2_X1 U658 ( .A1(n146), .A2(n98), .ZN(\ab[4][20] ) );
  NOR2_X1 U659 ( .A1(n137), .A2(n103), .ZN(\ab[6][18] ) );
  NOR2_X1 U660 ( .A1(n131), .A2(n110), .ZN(\ab[8][16] ) );
  NOR2_X1 U661 ( .A1(n127), .A2(n91), .ZN(\ab[10][14] ) );
  NOR2_X1 U662 ( .A1(n121), .A2(n64), .ZN(\ab[12][12] ) );
  NOR2_X1 U663 ( .A1(n115), .A2(n62), .ZN(\ab[14][10] ) );
  NOR2_X1 U664 ( .A1(n189), .A2(n60), .ZN(\ab[16][8] ) );
  NOR2_X1 U665 ( .A1(n182), .A2(n58), .ZN(\ab[18][6] ) );
  NOR2_X1 U666 ( .A1(n10), .A2(n55), .ZN(\ab[20][4] ) );
  NOR2_X1 U667 ( .A1(n123), .A2(n48), .ZN(\ab[27][13] ) );
  NOR2_X1 U668 ( .A1(n129), .A2(n50), .ZN(\ab[25][15] ) );
  NOR2_X1 U669 ( .A1(n135), .A2(n52), .ZN(\ab[23][17] ) );
  NOR2_X1 U670 ( .A1(n141), .A2(n54), .ZN(\ab[21][19] ) );
  NOR2_X1 U671 ( .A1(n151), .A2(n57), .ZN(\ab[19][21] ) );
  NOR2_X1 U672 ( .A1(n157), .A2(n59), .ZN(\ab[17][23] ) );
  NOR2_X1 U673 ( .A1(n162), .A2(n61), .ZN(\ab[15][25] ) );
  NOR2_X1 U674 ( .A1(n166), .A2(n63), .ZN(\ab[13][27] ) );
  NOR2_X1 U675 ( .A1(n170), .A2(n65), .ZN(\ab[11][29] ) );
  NOR2_X1 U676 ( .A1(n146), .A2(n96), .ZN(\ab[3][20] ) );
  NOR2_X1 U677 ( .A1(n137), .A2(n100), .ZN(\ab[5][18] ) );
  NOR2_X1 U678 ( .A1(n131), .A2(n107), .ZN(\ab[7][16] ) );
  NOR2_X1 U679 ( .A1(n195), .A2(n125), .ZN(\ab[9][14] ) );
  NOR2_X1 U680 ( .A1(n121), .A2(n65), .ZN(\ab[11][12] ) );
  NOR2_X1 U681 ( .A1(n115), .A2(n63), .ZN(\ab[13][10] ) );
  NOR2_X1 U682 ( .A1(n189), .A2(n61), .ZN(\ab[15][8] ) );
  NOR2_X1 U683 ( .A1(n126), .A2(n49), .ZN(\ab[26][14] ) );
  NOR2_X1 U684 ( .A1(n182), .A2(n59), .ZN(\ab[17][6] ) );
  NOR2_X1 U685 ( .A1(n132), .A2(n51), .ZN(\ab[24][16] ) );
  NOR2_X1 U686 ( .A1(n138), .A2(n53), .ZN(\ab[22][18] ) );
  NOR2_X1 U687 ( .A1(n147), .A2(n55), .ZN(\ab[20][20] ) );
  NOR2_X1 U688 ( .A1(n153), .A2(n58), .ZN(\ab[18][22] ) );
  NOR2_X1 U689 ( .A1(n158), .A2(n60), .ZN(\ab[16][24] ) );
  NOR2_X1 U690 ( .A1(n164), .A2(n62), .ZN(\ab[14][26] ) );
  NOR2_X1 U691 ( .A1(n168), .A2(n93), .ZN(\ab[12][28] ) );
  NOR2_X1 U692 ( .A1(n10), .A2(n57), .ZN(\ab[19][4] ) );
  NOR2_X1 U693 ( .A1(n137), .A2(n98), .ZN(\ab[4][18] ) );
  NOR2_X1 U694 ( .A1(n131), .A2(n104), .ZN(\ab[6][16] ) );
  NOR2_X1 U695 ( .A1(n125), .A2(n110), .ZN(\ab[8][14] ) );
  NOR2_X1 U696 ( .A1(n121), .A2(n91), .ZN(\ab[10][12] ) );
  NOR2_X1 U697 ( .A1(n115), .A2(n64), .ZN(\ab[12][10] ) );
  NOR2_X1 U698 ( .A1(n189), .A2(n62), .ZN(\ab[14][8] ) );
  NOR2_X1 U699 ( .A1(n183), .A2(n60), .ZN(\ab[16][6] ) );
  NOR2_X1 U700 ( .A1(n10), .A2(n58), .ZN(\ab[18][4] ) );
  NOR2_X1 U701 ( .A1(n137), .A2(n95), .ZN(\ab[3][18] ) );
  NOR2_X1 U702 ( .A1(n131), .A2(n101), .ZN(\ab[5][16] ) );
  NOR2_X1 U703 ( .A1(n125), .A2(n107), .ZN(\ab[7][14] ) );
  NOR2_X1 U704 ( .A1(n195), .A2(n119), .ZN(\ab[9][12] ) );
  NOR2_X1 U705 ( .A1(n115), .A2(n65), .ZN(\ab[11][10] ) );
  NOR2_X1 U706 ( .A1(n189), .A2(n63), .ZN(\ab[13][8] ) );
  NOR2_X1 U707 ( .A1(n183), .A2(n61), .ZN(\ab[15][6] ) );
  NOR2_X1 U708 ( .A1(n176), .A2(n59), .ZN(\ab[17][4] ) );
  NOR2_X1 U709 ( .A1(n129), .A2(n49), .ZN(\ab[26][15] ) );
  NOR2_X1 U710 ( .A1(n135), .A2(n51), .ZN(\ab[24][17] ) );
  NOR2_X1 U711 ( .A1(n141), .A2(n53), .ZN(\ab[22][19] ) );
  NOR2_X1 U712 ( .A1(n149), .A2(n55), .ZN(\ab[20][21] ) );
  NOR2_X1 U713 ( .A1(n155), .A2(n58), .ZN(\ab[18][23] ) );
  NOR2_X1 U714 ( .A1(n161), .A2(n60), .ZN(\ab[16][25] ) );
  NOR2_X1 U715 ( .A1(n166), .A2(n62), .ZN(\ab[14][27] ) );
  NOR2_X1 U716 ( .A1(n170), .A2(n93), .ZN(\ab[12][29] ) );
  NOR2_X1 U717 ( .A1(n126), .A2(n48), .ZN(\ab[27][14] ) );
  NOR2_X1 U718 ( .A1(n132), .A2(n50), .ZN(\ab[25][16] ) );
  NOR2_X1 U719 ( .A1(n138), .A2(n52), .ZN(\ab[23][18] ) );
  NOR2_X1 U720 ( .A1(n147), .A2(n54), .ZN(\ab[21][20] ) );
  NOR2_X1 U721 ( .A1(n153), .A2(n57), .ZN(\ab[19][22] ) );
  NOR2_X1 U722 ( .A1(n158), .A2(n59), .ZN(\ab[17][24] ) );
  NOR2_X1 U723 ( .A1(n163), .A2(n61), .ZN(\ab[15][26] ) );
  NOR2_X1 U724 ( .A1(n169), .A2(n63), .ZN(\ab[13][28] ) );
  NOR2_X1 U725 ( .A1(n125), .A2(n47), .ZN(\ab[28][14] ) );
  NOR2_X1 U726 ( .A1(n132), .A2(n49), .ZN(\ab[26][16] ) );
  NOR2_X1 U727 ( .A1(n138), .A2(n51), .ZN(\ab[24][18] ) );
  NOR2_X1 U728 ( .A1(n147), .A2(n53), .ZN(\ab[22][20] ) );
  NOR2_X1 U729 ( .A1(n153), .A2(n55), .ZN(\ab[20][22] ) );
  NOR2_X1 U730 ( .A1(n160), .A2(n58), .ZN(\ab[18][24] ) );
  NOR2_X1 U731 ( .A1(n163), .A2(n60), .ZN(\ab[16][26] ) );
  NOR2_X1 U732 ( .A1(n169), .A2(n62), .ZN(\ab[14][28] ) );
  NOR2_X1 U733 ( .A1(n129), .A2(n48), .ZN(\ab[27][15] ) );
  NOR2_X1 U734 ( .A1(n135), .A2(n50), .ZN(\ab[25][17] ) );
  NOR2_X1 U735 ( .A1(n141), .A2(n52), .ZN(\ab[23][19] ) );
  NOR2_X1 U736 ( .A1(n150), .A2(n54), .ZN(\ab[21][21] ) );
  NOR2_X1 U737 ( .A1(n157), .A2(n57), .ZN(\ab[19][23] ) );
  NOR2_X1 U738 ( .A1(n162), .A2(n59), .ZN(\ab[17][25] ) );
  NOR2_X1 U739 ( .A1(n166), .A2(n61), .ZN(\ab[15][27] ) );
  NOR2_X1 U740 ( .A1(n170), .A2(n63), .ZN(\ab[13][29] ) );
  NOR2_X1 U741 ( .A1(n131), .A2(n98), .ZN(\ab[4][16] ) );
  NOR2_X1 U742 ( .A1(n125), .A2(n104), .ZN(\ab[6][14] ) );
  NOR2_X1 U743 ( .A1(n119), .A2(n110), .ZN(\ab[8][12] ) );
  NOR2_X1 U744 ( .A1(n115), .A2(n91), .ZN(\ab[10][10] ) );
  NOR2_X1 U745 ( .A1(n189), .A2(n93), .ZN(\ab[12][8] ) );
  NOR2_X1 U746 ( .A1(n183), .A2(n62), .ZN(\ab[14][6] ) );
  NOR2_X1 U747 ( .A1(n177), .A2(n60), .ZN(\ab[16][4] ) );
  NOR2_X1 U748 ( .A1(n131), .A2(n96), .ZN(\ab[3][16] ) );
  NOR2_X1 U749 ( .A1(n125), .A2(n101), .ZN(\ab[5][14] ) );
  NOR2_X1 U750 ( .A1(n119), .A2(n107), .ZN(\ab[7][12] ) );
  NOR2_X1 U751 ( .A1(n128), .A2(n47), .ZN(\ab[28][15] ) );
  NOR2_X1 U752 ( .A1(n195), .A2(n113), .ZN(\ab[9][10] ) );
  NOR2_X1 U753 ( .A1(n135), .A2(n49), .ZN(\ab[26][17] ) );
  NOR2_X1 U754 ( .A1(n189), .A2(n65), .ZN(\ab[11][8] ) );
  NOR2_X1 U755 ( .A1(n141), .A2(n51), .ZN(\ab[24][19] ) );
  NOR2_X1 U756 ( .A1(n183), .A2(n63), .ZN(\ab[13][6] ) );
  NOR2_X1 U757 ( .A1(n151), .A2(n53), .ZN(\ab[22][21] ) );
  NOR2_X1 U758 ( .A1(n155), .A2(n55), .ZN(\ab[20][23] ) );
  NOR2_X1 U759 ( .A1(n162), .A2(n58), .ZN(\ab[18][25] ) );
  NOR2_X1 U760 ( .A1(n167), .A2(n60), .ZN(\ab[16][27] ) );
  NOR2_X1 U761 ( .A1(n170), .A2(n62), .ZN(\ab[14][29] ) );
  NOR2_X1 U762 ( .A1(n177), .A2(n61), .ZN(\ab[15][4] ) );
  NOR2_X1 U763 ( .A1(n132), .A2(n48), .ZN(\ab[27][16] ) );
  NOR2_X1 U764 ( .A1(n138), .A2(n50), .ZN(\ab[25][18] ) );
  NOR2_X1 U765 ( .A1(n147), .A2(n52), .ZN(\ab[23][20] ) );
  NOR2_X1 U766 ( .A1(n153), .A2(n54), .ZN(\ab[21][22] ) );
  NOR2_X1 U767 ( .A1(n158), .A2(n57), .ZN(\ab[19][24] ) );
  NOR2_X1 U768 ( .A1(n163), .A2(n59), .ZN(\ab[17][26] ) );
  NOR2_X1 U769 ( .A1(n169), .A2(n61), .ZN(\ab[15][28] ) );
  NOR2_X1 U770 ( .A1(n125), .A2(n98), .ZN(\ab[4][14] ) );
  NOR2_X1 U771 ( .A1(n119), .A2(n104), .ZN(\ab[6][12] ) );
  NOR2_X1 U772 ( .A1(n113), .A2(n110), .ZN(\ab[8][10] ) );
  NOR2_X1 U773 ( .A1(n189), .A2(n89), .ZN(\ab[10][8] ) );
  NOR2_X1 U774 ( .A1(n183), .A2(n93), .ZN(\ab[12][6] ) );
  NOR2_X1 U775 ( .A1(n177), .A2(n62), .ZN(\ab[14][4] ) );
  NOR2_X1 U776 ( .A1(n125), .A2(n95), .ZN(\ab[3][14] ) );
  NOR2_X1 U777 ( .A1(n119), .A2(n101), .ZN(\ab[5][12] ) );
  NOR2_X1 U778 ( .A1(n113), .A2(n107), .ZN(\ab[7][10] ) );
  NOR2_X1 U779 ( .A1(n193), .A2(n187), .ZN(\ab[9][8] ) );
  NOR2_X1 U780 ( .A1(n183), .A2(n65), .ZN(\ab[11][6] ) );
  NOR2_X1 U781 ( .A1(n177), .A2(n63), .ZN(\ab[13][4] ) );
  NOR2_X1 U782 ( .A1(n131), .A2(n47), .ZN(\ab[28][16] ) );
  NOR2_X1 U783 ( .A1(n138), .A2(n49), .ZN(\ab[26][18] ) );
  NOR2_X1 U784 ( .A1(n147), .A2(n51), .ZN(\ab[24][20] ) );
  NOR2_X1 U785 ( .A1(n153), .A2(n53), .ZN(\ab[22][22] ) );
  NOR2_X1 U786 ( .A1(n158), .A2(n55), .ZN(\ab[20][24] ) );
  NOR2_X1 U787 ( .A1(n164), .A2(n58), .ZN(\ab[18][26] ) );
  NOR2_X1 U788 ( .A1(n169), .A2(n60), .ZN(\ab[16][28] ) );
  NOR2_X1 U789 ( .A1(n119), .A2(n98), .ZN(\ab[4][12] ) );
  NOR2_X1 U790 ( .A1(n113), .A2(n104), .ZN(\ab[6][10] ) );
  NOR2_X1 U791 ( .A1(n187), .A2(n108), .ZN(\ab[8][8] ) );
  NOR2_X1 U792 ( .A1(n183), .A2(n89), .ZN(\ab[10][6] ) );
  NOR2_X1 U793 ( .A1(n177), .A2(n93), .ZN(\ab[12][4] ) );
  NOR2_X1 U794 ( .A1(n135), .A2(n48), .ZN(\ab[27][17] ) );
  NOR2_X1 U795 ( .A1(n141), .A2(n50), .ZN(\ab[25][19] ) );
  NOR2_X1 U796 ( .A1(n149), .A2(n52), .ZN(\ab[23][21] ) );
  NOR2_X1 U797 ( .A1(n157), .A2(n54), .ZN(\ab[21][23] ) );
  NOR2_X1 U798 ( .A1(n161), .A2(n57), .ZN(\ab[19][25] ) );
  NOR2_X1 U799 ( .A1(n166), .A2(n59), .ZN(\ab[17][27] ) );
  NOR2_X1 U800 ( .A1(n170), .A2(n61), .ZN(\ab[15][29] ) );
  NOR2_X1 U801 ( .A1(n131), .A2(n46), .ZN(\ab[29][16] ) );
  NOR2_X1 U802 ( .A1(n119), .A2(n95), .ZN(\ab[3][12] ) );
  NOR2_X1 U803 ( .A1(n113), .A2(n101), .ZN(\ab[5][10] ) );
  NOR2_X1 U804 ( .A1(n187), .A2(n105), .ZN(\ab[7][8] ) );
  NOR2_X1 U805 ( .A1(n193), .A2(n181), .ZN(\ab[9][6] ) );
  NOR2_X1 U806 ( .A1(n177), .A2(n65), .ZN(\ab[11][4] ) );
  NOR2_X1 U807 ( .A1(n113), .A2(n98), .ZN(\ab[4][10] ) );
  NOR2_X1 U808 ( .A1(n187), .A2(n102), .ZN(\ab[6][8] ) );
  NOR2_X1 U809 ( .A1(n181), .A2(n108), .ZN(\ab[8][6] ) );
  NOR2_X1 U810 ( .A1(n177), .A2(n89), .ZN(\ab[10][4] ) );
  NOR2_X1 U811 ( .A1(n113), .A2(n96), .ZN(\ab[3][10] ) );
  NOR2_X1 U812 ( .A1(n187), .A2(n99), .ZN(\ab[5][8] ) );
  NOR2_X1 U813 ( .A1(n181), .A2(n105), .ZN(\ab[7][6] ) );
  NOR2_X1 U814 ( .A1(n193), .A2(n176), .ZN(\ab[9][4] ) );
  NOR2_X1 U815 ( .A1(n187), .A2(n97), .ZN(\ab[4][8] ) );
  NOR2_X1 U816 ( .A1(n181), .A2(n102), .ZN(\ab[6][6] ) );
  NOR2_X1 U817 ( .A1(n176), .A2(n108), .ZN(\ab[8][4] ) );
  NOR2_X1 U818 ( .A1(n187), .A2(n96), .ZN(\ab[3][8] ) );
  NOR2_X1 U819 ( .A1(n181), .A2(n99), .ZN(\ab[5][6] ) );
  NOR2_X1 U820 ( .A1(n176), .A2(n105), .ZN(\ab[7][4] ) );
  NOR2_X1 U821 ( .A1(n134), .A2(n47), .ZN(\ab[28][17] ) );
  NOR2_X1 U822 ( .A1(n141), .A2(n49), .ZN(\ab[26][19] ) );
  NOR2_X1 U823 ( .A1(n150), .A2(n51), .ZN(\ab[24][21] ) );
  NOR2_X1 U824 ( .A1(n155), .A2(n53), .ZN(\ab[22][23] ) );
  NOR2_X1 U825 ( .A1(n162), .A2(n55), .ZN(\ab[20][25] ) );
  NOR2_X1 U826 ( .A1(n167), .A2(n58), .ZN(\ab[18][27] ) );
  NOR2_X1 U827 ( .A1(n170), .A2(n60), .ZN(\ab[16][29] ) );
  NOR2_X1 U828 ( .A1(n138), .A2(n48), .ZN(\ab[27][18] ) );
  NOR2_X1 U829 ( .A1(n147), .A2(n50), .ZN(\ab[25][20] ) );
  NOR2_X1 U830 ( .A1(n153), .A2(n52), .ZN(\ab[23][22] ) );
  NOR2_X1 U831 ( .A1(n160), .A2(n54), .ZN(\ab[21][24] ) );
  NOR2_X1 U832 ( .A1(n163), .A2(n57), .ZN(\ab[19][26] ) );
  NOR2_X1 U833 ( .A1(n168), .A2(n59), .ZN(\ab[17][28] ) );
  NOR2_X1 U834 ( .A1(n181), .A2(n97), .ZN(\ab[4][6] ) );
  NOR2_X1 U835 ( .A1(n176), .A2(n102), .ZN(\ab[6][4] ) );
  NOR2_X1 U836 ( .A1(n181), .A2(n95), .ZN(\ab[3][6] ) );
  NOR2_X1 U837 ( .A1(n176), .A2(n99), .ZN(\ab[5][4] ) );
  NOR2_X1 U838 ( .A1(n176), .A2(n97), .ZN(\ab[4][4] ) );
  NOR2_X1 U839 ( .A1(n176), .A2(n95), .ZN(\ab[3][4] ) );
  NOR2_X1 U840 ( .A1(n134), .A2(n46), .ZN(\ab[29][17] ) );
  NOR2_X1 U841 ( .A1(n137), .A2(n47), .ZN(\ab[28][18] ) );
  NOR2_X1 U842 ( .A1(n147), .A2(n49), .ZN(\ab[26][20] ) );
  NOR2_X1 U843 ( .A1(n153), .A2(n51), .ZN(\ab[24][22] ) );
  NOR2_X1 U844 ( .A1(n158), .A2(n53), .ZN(\ab[22][24] ) );
  NOR2_X1 U845 ( .A1(n163), .A2(n55), .ZN(\ab[20][26] ) );
  NOR2_X1 U846 ( .A1(n169), .A2(n58), .ZN(\ab[18][28] ) );
  NOR2_X1 U847 ( .A1(n141), .A2(n48), .ZN(\ab[27][19] ) );
  NOR2_X1 U848 ( .A1(n151), .A2(n50), .ZN(\ab[25][21] ) );
  NOR2_X1 U849 ( .A1(n157), .A2(n52), .ZN(\ab[23][23] ) );
  NOR2_X1 U850 ( .A1(n162), .A2(n54), .ZN(\ab[21][25] ) );
  NOR2_X1 U851 ( .A1(n166), .A2(n57), .ZN(\ab[19][27] ) );
  NOR2_X1 U852 ( .A1(n170), .A2(n59), .ZN(\ab[17][29] ) );
  NOR2_X1 U853 ( .A1(n137), .A2(n46), .ZN(\ab[29][18] ) );
  NOR2_X1 U854 ( .A1(n140), .A2(n47), .ZN(\ab[28][19] ) );
  NOR2_X1 U855 ( .A1(n149), .A2(n49), .ZN(\ab[26][21] ) );
  NOR2_X1 U856 ( .A1(n155), .A2(n51), .ZN(\ab[24][23] ) );
  NOR2_X1 U857 ( .A1(n161), .A2(n53), .ZN(\ab[22][25] ) );
  NOR2_X1 U858 ( .A1(n167), .A2(n55), .ZN(\ab[20][27] ) );
  NOR2_X1 U859 ( .A1(n170), .A2(n58), .ZN(\ab[18][29] ) );
  NOR2_X1 U860 ( .A1(n147), .A2(n48), .ZN(\ab[27][20] ) );
  NOR2_X1 U861 ( .A1(n153), .A2(n50), .ZN(\ab[25][22] ) );
  NOR2_X1 U862 ( .A1(n160), .A2(n52), .ZN(\ab[23][24] ) );
  NOR2_X1 U863 ( .A1(n164), .A2(n54), .ZN(\ab[21][26] ) );
  NOR2_X1 U864 ( .A1(n168), .A2(n57), .ZN(\ab[19][28] ) );
  NOR2_X1 U865 ( .A1(n173), .A2(n44), .ZN(\ab[30][3] ) );
  NOR2_X1 U866 ( .A1(n178), .A2(n44), .ZN(\ab[30][5] ) );
  NOR2_X1 U867 ( .A1(n116), .A2(n44), .ZN(\ab[30][11] ) );
  NOR2_X1 U868 ( .A1(n171), .A2(n44), .ZN(\ab[30][2] ) );
  NOR2_X1 U869 ( .A1(n190), .A2(n46), .ZN(\ab[29][9] ) );
  NOR2_X1 U870 ( .A1(n173), .A2(n46), .ZN(\ab[29][3] ) );
  NOR2_X1 U871 ( .A1(n143), .A2(n44), .ZN(\ab[30][1] ) );
  NOR2_X1 U872 ( .A1(n171), .A2(n46), .ZN(\ab[29][2] ) );
  NOR2_X1 U873 ( .A1(n173), .A2(n47), .ZN(\ab[28][3] ) );
  NOR2_X1 U874 ( .A1(n155), .A2(n109), .ZN(\ab[8][23] ) );
  NOR2_X1 U875 ( .A1(n194), .A2(n157), .ZN(\ab[9][23] ) );
  NOR2_X1 U876 ( .A1(n151), .A2(n90), .ZN(\ab[10][21] ) );
  NOR2_X1 U877 ( .A1(n149), .A2(n92), .ZN(\ab[11][21] ) );
  NOR2_X1 U878 ( .A1(n142), .A2(n64), .ZN(\ab[12][19] ) );
  NOR2_X1 U879 ( .A1(n142), .A2(n63), .ZN(\ab[13][19] ) );
  NOR2_X1 U880 ( .A1(n136), .A2(n62), .ZN(\ab[14][17] ) );
  NOR2_X1 U881 ( .A1(n136), .A2(n61), .ZN(\ab[15][17] ) );
  NOR2_X1 U882 ( .A1(n130), .A2(n60), .ZN(\ab[16][15] ) );
  NOR2_X1 U883 ( .A1(n129), .A2(n59), .ZN(\ab[17][15] ) );
  NOR2_X1 U884 ( .A1(n123), .A2(n58), .ZN(\ab[18][13] ) );
  NOR2_X1 U885 ( .A1(n123), .A2(n57), .ZN(\ab[19][13] ) );
  NOR2_X1 U886 ( .A1(n117), .A2(n55), .ZN(\ab[20][11] ) );
  NOR2_X1 U887 ( .A1(n117), .A2(n54), .ZN(\ab[21][11] ) );
  NOR2_X1 U888 ( .A1(n191), .A2(n53), .ZN(\ab[22][9] ) );
  NOR2_X1 U889 ( .A1(n191), .A2(n52), .ZN(\ab[23][9] ) );
  NOR2_X1 U890 ( .A1(n185), .A2(n51), .ZN(\ab[24][7] ) );
  NOR2_X1 U891 ( .A1(n179), .A2(n48), .ZN(\ab[27][5] ) );
  NOR2_X1 U892 ( .A1(n179), .A2(n49), .ZN(\ab[26][5] ) );
  NOR2_X1 U893 ( .A1(n155), .A2(n103), .ZN(\ab[6][23] ) );
  NOR2_X1 U894 ( .A1(n149), .A2(n109), .ZN(\ab[8][21] ) );
  NOR2_X1 U895 ( .A1(n194), .A2(n150), .ZN(\ab[9][21] ) );
  NOR2_X1 U896 ( .A1(n142), .A2(n90), .ZN(\ab[10][19] ) );
  NOR2_X1 U897 ( .A1(n142), .A2(n92), .ZN(\ab[11][19] ) );
  NOR2_X1 U898 ( .A1(n136), .A2(n64), .ZN(\ab[12][17] ) );
  NOR2_X1 U899 ( .A1(n136), .A2(n63), .ZN(\ab[13][17] ) );
  NOR2_X1 U900 ( .A1(n130), .A2(n62), .ZN(\ab[14][15] ) );
  NOR2_X1 U901 ( .A1(n130), .A2(n61), .ZN(\ab[15][15] ) );
  NOR2_X1 U902 ( .A1(n124), .A2(n60), .ZN(\ab[16][13] ) );
  NOR2_X1 U903 ( .A1(n123), .A2(n59), .ZN(\ab[17][13] ) );
  NOR2_X1 U904 ( .A1(n117), .A2(n57), .ZN(\ab[19][11] ) );
  NOR2_X1 U905 ( .A1(n117), .A2(n58), .ZN(\ab[18][11] ) );
  NOR2_X1 U906 ( .A1(n191), .A2(n54), .ZN(\ab[21][9] ) );
  NOR2_X1 U907 ( .A1(n191), .A2(n55), .ZN(\ab[20][9] ) );
  NOR2_X1 U908 ( .A1(n185), .A2(n52), .ZN(\ab[23][7] ) );
  NOR2_X1 U909 ( .A1(n185), .A2(n53), .ZN(\ab[22][7] ) );
  NOR2_X1 U910 ( .A1(n179), .A2(n50), .ZN(\ab[25][5] ) );
  NOR2_X1 U911 ( .A1(n179), .A2(n51), .ZN(\ab[24][5] ) );
  NOR2_X1 U912 ( .A1(n162), .A2(n95), .ZN(\ab[3][25] ) );
  NOR2_X1 U913 ( .A1(n157), .A2(n100), .ZN(\ab[5][23] ) );
  NOR2_X1 U914 ( .A1(n151), .A2(n106), .ZN(\ab[7][21] ) );
  NOR2_X1 U915 ( .A1(n194), .A2(n140), .ZN(\ab[9][19] ) );
  NOR2_X1 U916 ( .A1(n136), .A2(n92), .ZN(\ab[11][17] ) );
  NOR2_X1 U917 ( .A1(n130), .A2(n63), .ZN(\ab[13][15] ) );
  NOR2_X1 U918 ( .A1(n124), .A2(n61), .ZN(\ab[15][13] ) );
  NOR2_X1 U919 ( .A1(n117), .A2(n59), .ZN(\ab[17][11] ) );
  NOR2_X1 U920 ( .A1(n191), .A2(n57), .ZN(\ab[19][9] ) );
  NOR2_X1 U921 ( .A1(n185), .A2(n54), .ZN(\ab[21][7] ) );
  NOR2_X1 U922 ( .A1(n179), .A2(n52), .ZN(\ab[23][5] ) );
  NOR2_X1 U923 ( .A1(n174), .A2(n48), .ZN(\ab[27][3] ) );
  NOR2_X1 U924 ( .A1(n174), .A2(n49), .ZN(\ab[26][3] ) );
  NOR2_X1 U925 ( .A1(n155), .A2(n98), .ZN(\ab[4][23] ) );
  NOR2_X1 U926 ( .A1(n150), .A2(n103), .ZN(\ab[6][21] ) );
  NOR2_X1 U927 ( .A1(n140), .A2(n109), .ZN(\ab[8][19] ) );
  NOR2_X1 U928 ( .A1(n136), .A2(n90), .ZN(\ab[10][17] ) );
  NOR2_X1 U929 ( .A1(n130), .A2(n93), .ZN(\ab[12][15] ) );
  NOR2_X1 U930 ( .A1(n124), .A2(n62), .ZN(\ab[14][13] ) );
  NOR2_X1 U931 ( .A1(n118), .A2(n60), .ZN(\ab[16][11] ) );
  NOR2_X1 U932 ( .A1(n191), .A2(n58), .ZN(\ab[18][9] ) );
  NOR2_X1 U933 ( .A1(n185), .A2(n55), .ZN(\ab[20][7] ) );
  NOR2_X1 U934 ( .A1(n179), .A2(n53), .ZN(\ab[22][5] ) );
  NOR2_X1 U935 ( .A1(n174), .A2(n50), .ZN(\ab[25][3] ) );
  NOR2_X1 U936 ( .A1(n174), .A2(n51), .ZN(\ab[24][3] ) );
  NOR2_X1 U937 ( .A1(n171), .A2(n47), .ZN(\ab[28][2] ) );
  NOR2_X1 U938 ( .A1(n157), .A2(n96), .ZN(\ab[3][23] ) );
  NOR2_X1 U939 ( .A1(n140), .A2(n106), .ZN(\ab[7][19] ) );
  NOR2_X1 U940 ( .A1(n194), .A2(n134), .ZN(\ab[9][17] ) );
  NOR2_X1 U941 ( .A1(n130), .A2(n65), .ZN(\ab[11][15] ) );
  NOR2_X1 U942 ( .A1(n124), .A2(n63), .ZN(\ab[13][13] ) );
  NOR2_X1 U943 ( .A1(n118), .A2(n61), .ZN(\ab[15][11] ) );
  NOR2_X1 U944 ( .A1(n191), .A2(n59), .ZN(\ab[17][9] ) );
  NOR2_X1 U945 ( .A1(n185), .A2(n57), .ZN(\ab[19][7] ) );
  NOR2_X1 U946 ( .A1(n179), .A2(n54), .ZN(\ab[21][5] ) );
  NOR2_X1 U947 ( .A1(n14), .A2(n48), .ZN(\ab[27][2] ) );
  NOR2_X1 U948 ( .A1(n14), .A2(n49), .ZN(\ab[26][2] ) );
  NOR2_X1 U949 ( .A1(n151), .A2(n98), .ZN(\ab[4][21] ) );
  NOR2_X1 U950 ( .A1(n140), .A2(n103), .ZN(\ab[6][19] ) );
  NOR2_X1 U951 ( .A1(n134), .A2(n109), .ZN(\ab[8][17] ) );
  NOR2_X1 U952 ( .A1(n130), .A2(n91), .ZN(\ab[10][15] ) );
  NOR2_X1 U953 ( .A1(n124), .A2(n64), .ZN(\ab[12][13] ) );
  NOR2_X1 U954 ( .A1(n118), .A2(n62), .ZN(\ab[14][11] ) );
  NOR2_X1 U955 ( .A1(n192), .A2(n60), .ZN(\ab[16][9] ) );
  NOR2_X1 U956 ( .A1(n185), .A2(n58), .ZN(\ab[18][7] ) );
  NOR2_X1 U957 ( .A1(n179), .A2(n55), .ZN(\ab[20][5] ) );
  NOR2_X1 U958 ( .A1(n174), .A2(n52), .ZN(\ab[23][3] ) );
  NOR2_X1 U959 ( .A1(n14), .A2(n50), .ZN(\ab[25][2] ) );
  NOR2_X1 U960 ( .A1(n174), .A2(n53), .ZN(\ab[22][3] ) );
  NOR2_X1 U961 ( .A1(n150), .A2(n96), .ZN(\ab[3][21] ) );
  NOR2_X1 U962 ( .A1(n140), .A2(n100), .ZN(\ab[5][19] ) );
  NOR2_X1 U963 ( .A1(n134), .A2(n106), .ZN(\ab[7][17] ) );
  NOR2_X1 U964 ( .A1(n195), .A2(n128), .ZN(\ab[9][15] ) );
  NOR2_X1 U965 ( .A1(n124), .A2(n65), .ZN(\ab[11][13] ) );
  NOR2_X1 U966 ( .A1(n118), .A2(n63), .ZN(\ab[13][11] ) );
  NOR2_X1 U967 ( .A1(n192), .A2(n61), .ZN(\ab[15][9] ) );
  NOR2_X1 U968 ( .A1(n185), .A2(n59), .ZN(\ab[17][7] ) );
  NOR2_X1 U969 ( .A1(n179), .A2(n57), .ZN(\ab[19][5] ) );
  NOR2_X1 U970 ( .A1(n143), .A2(n46), .ZN(\ab[29][1] ) );
  NOR2_X1 U971 ( .A1(n149), .A2(net144909), .ZN(\ab[2][21] ) );
  AND2_X1 U972 ( .A1(\ab[1][21] ), .A2(\ab[0][22] ), .ZN(\CARRYB[1][21] ) );
  NOR2_X1 U973 ( .A1(n140), .A2(n98), .ZN(\ab[4][19] ) );
  NOR2_X1 U974 ( .A1(n134), .A2(n103), .ZN(\ab[6][17] ) );
  NOR2_X1 U975 ( .A1(n128), .A2(n110), .ZN(\ab[8][15] ) );
  NOR2_X1 U976 ( .A1(n124), .A2(n91), .ZN(\ab[10][13] ) );
  NOR2_X1 U977 ( .A1(n118), .A2(n64), .ZN(\ab[12][11] ) );
  NOR2_X1 U978 ( .A1(n192), .A2(n62), .ZN(\ab[14][9] ) );
  NOR2_X1 U979 ( .A1(n186), .A2(n60), .ZN(\ab[16][7] ) );
  NOR2_X1 U980 ( .A1(n179), .A2(n58), .ZN(\ab[18][5] ) );
  NOR2_X1 U981 ( .A1(n174), .A2(n54), .ZN(\ab[21][3] ) );
  NOR2_X1 U982 ( .A1(n14), .A2(n51), .ZN(\ab[24][2] ) );
  NOR2_X1 U983 ( .A1(n140), .A2(n96), .ZN(\ab[3][19] ) );
  NOR2_X1 U984 ( .A1(n134), .A2(n100), .ZN(\ab[5][17] ) );
  NOR2_X1 U985 ( .A1(n128), .A2(n107), .ZN(\ab[7][15] ) );
  NOR2_X1 U986 ( .A1(n195), .A2(n122), .ZN(\ab[9][13] ) );
  NOR2_X1 U987 ( .A1(n118), .A2(n65), .ZN(\ab[11][11] ) );
  NOR2_X1 U988 ( .A1(n192), .A2(n63), .ZN(\ab[13][9] ) );
  NOR2_X1 U989 ( .A1(n186), .A2(n61), .ZN(\ab[15][7] ) );
  NOR2_X1 U990 ( .A1(n179), .A2(n59), .ZN(\ab[17][5] ) );
  NOR2_X1 U991 ( .A1(n140), .A2(net144909), .ZN(\ab[2][19] ) );
  AND2_X1 U992 ( .A1(\ab[1][19] ), .A2(\ab[0][20] ), .ZN(\CARRYB[1][19] ) );
  NOR2_X1 U993 ( .A1(n134), .A2(n98), .ZN(\ab[4][17] ) );
  NOR2_X1 U994 ( .A1(n128), .A2(n104), .ZN(\ab[6][15] ) );
  NOR2_X1 U995 ( .A1(n122), .A2(n110), .ZN(\ab[8][13] ) );
  NOR2_X1 U996 ( .A1(n118), .A2(n91), .ZN(\ab[10][11] ) );
  NOR2_X1 U997 ( .A1(n192), .A2(n93), .ZN(\ab[12][9] ) );
  NOR2_X1 U998 ( .A1(n186), .A2(n62), .ZN(\ab[14][7] ) );
  NOR2_X1 U999 ( .A1(n180), .A2(n60), .ZN(\ab[16][5] ) );
  NOR2_X1 U1000 ( .A1(n174), .A2(n55), .ZN(\ab[20][3] ) );
  NOR2_X1 U1001 ( .A1(n14), .A2(n52), .ZN(\ab[23][2] ) );
  NOR2_X1 U1002 ( .A1(n174), .A2(n57), .ZN(\ab[19][3] ) );
  NOR2_X1 U1003 ( .A1(n143), .A2(n47), .ZN(\ab[28][1] ) );
  NOR2_X1 U1004 ( .A1(n14), .A2(n53), .ZN(\ab[22][2] ) );
  NOR2_X1 U1005 ( .A1(n144), .A2(n48), .ZN(\ab[27][1] ) );
  NOR2_X1 U1006 ( .A1(n174), .A2(n58), .ZN(\ab[18][3] ) );
  NOR2_X1 U1007 ( .A1(n14), .A2(n54), .ZN(\ab[21][2] ) );
  NOR2_X1 U1008 ( .A1(n144), .A2(n49), .ZN(\ab[26][1] ) );
  NOR2_X1 U1009 ( .A1(n14), .A2(n55), .ZN(\ab[20][2] ) );
  NOR2_X1 U1010 ( .A1(n134), .A2(n95), .ZN(\ab[3][17] ) );
  NOR2_X1 U1011 ( .A1(n128), .A2(n101), .ZN(\ab[5][15] ) );
  NOR2_X1 U1012 ( .A1(n122), .A2(n107), .ZN(\ab[7][13] ) );
  NOR2_X1 U1013 ( .A1(n195), .A2(n116), .ZN(\ab[9][11] ) );
  NOR2_X1 U1014 ( .A1(n192), .A2(n65), .ZN(\ab[11][9] ) );
  NOR2_X1 U1015 ( .A1(n186), .A2(n63), .ZN(\ab[13][7] ) );
  NOR2_X1 U1016 ( .A1(n180), .A2(n61), .ZN(\ab[15][5] ) );
  NOR2_X1 U1017 ( .A1(n134), .A2(net144909), .ZN(\ab[2][17] ) );
  AND2_X1 U1018 ( .A1(\ab[1][17] ), .A2(\ab[0][18] ), .ZN(\CARRYB[1][17] ) );
  NOR2_X1 U1019 ( .A1(n128), .A2(n98), .ZN(\ab[4][15] ) );
  NOR2_X1 U1020 ( .A1(n122), .A2(n104), .ZN(\ab[6][13] ) );
  NOR2_X1 U1021 ( .A1(n116), .A2(n110), .ZN(\ab[8][11] ) );
  NOR2_X1 U1022 ( .A1(n192), .A2(n89), .ZN(\ab[10][9] ) );
  NOR2_X1 U1023 ( .A1(n186), .A2(n93), .ZN(\ab[12][7] ) );
  NOR2_X1 U1024 ( .A1(n180), .A2(n62), .ZN(\ab[14][5] ) );
  NOR2_X1 U1025 ( .A1(n172), .A2(n57), .ZN(\ab[19][2] ) );
  NOR2_X1 U1026 ( .A1(n174), .A2(n59), .ZN(\ab[17][3] ) );
  NOR2_X1 U1027 ( .A1(n144), .A2(n50), .ZN(\ab[25][1] ) );
  NOR2_X1 U1028 ( .A1(n144), .A2(n51), .ZN(\ab[24][1] ) );
  NOR2_X1 U1029 ( .A1(n175), .A2(n60), .ZN(\ab[16][3] ) );
  NOR2_X1 U1030 ( .A1(n128), .A2(n95), .ZN(\ab[3][15] ) );
  NOR2_X1 U1031 ( .A1(n122), .A2(n101), .ZN(\ab[5][13] ) );
  NOR2_X1 U1032 ( .A1(n116), .A2(n107), .ZN(\ab[7][11] ) );
  NOR2_X1 U1033 ( .A1(n193), .A2(n190), .ZN(\ab[9][9] ) );
  NOR2_X1 U1034 ( .A1(n186), .A2(n65), .ZN(\ab[11][7] ) );
  NOR2_X1 U1035 ( .A1(n180), .A2(n63), .ZN(\ab[13][5] ) );
  NOR2_X1 U1036 ( .A1(n128), .A2(net144909), .ZN(\ab[2][15] ) );
  AND2_X1 U1037 ( .A1(\ab[1][15] ), .A2(\ab[0][16] ), .ZN(\CARRYB[1][15] ) );
  NOR2_X1 U1038 ( .A1(n122), .A2(n98), .ZN(\ab[4][13] ) );
  NOR2_X1 U1039 ( .A1(n116), .A2(n104), .ZN(\ab[6][11] ) );
  NOR2_X1 U1040 ( .A1(n190), .A2(n108), .ZN(\ab[8][9] ) );
  NOR2_X1 U1041 ( .A1(n186), .A2(n89), .ZN(\ab[10][7] ) );
  NOR2_X1 U1042 ( .A1(n180), .A2(n93), .ZN(\ab[12][5] ) );
  NOR2_X1 U1043 ( .A1(n144), .A2(n52), .ZN(\ab[23][1] ) );
  NOR2_X1 U1044 ( .A1(n175), .A2(n61), .ZN(\ab[15][3] ) );
  NOR2_X1 U1045 ( .A1(n172), .A2(n58), .ZN(\ab[18][2] ) );
  NOR2_X1 U1046 ( .A1(n144), .A2(n53), .ZN(\ab[22][1] ) );
  NOR2_X1 U1047 ( .A1(n172), .A2(n59), .ZN(\ab[17][2] ) );
  NOR2_X1 U1048 ( .A1(n175), .A2(n62), .ZN(\ab[14][3] ) );
  NOR2_X1 U1049 ( .A1(n144), .A2(n54), .ZN(\ab[21][1] ) );
  NOR2_X1 U1050 ( .A1(n122), .A2(n96), .ZN(\ab[3][13] ) );
  NOR2_X1 U1051 ( .A1(n116), .A2(n101), .ZN(\ab[5][11] ) );
  NOR2_X1 U1052 ( .A1(n190), .A2(n105), .ZN(\ab[7][9] ) );
  NOR2_X1 U1053 ( .A1(n193), .A2(n184), .ZN(\ab[9][7] ) );
  NOR2_X1 U1054 ( .A1(n180), .A2(n65), .ZN(\ab[11][5] ) );
  NOR2_X1 U1055 ( .A1(n172), .A2(n60), .ZN(\ab[16][2] ) );
  NOR2_X1 U1056 ( .A1(n144), .A2(n55), .ZN(\ab[20][1] ) );
  NOR2_X1 U1057 ( .A1(n175), .A2(n63), .ZN(\ab[13][3] ) );
  NOR2_X1 U1058 ( .A1(n122), .A2(net144909), .ZN(\ab[2][13] ) );
  AND2_X1 U1059 ( .A1(\ab[1][13] ), .A2(\ab[0][14] ), .ZN(\CARRYB[1][13] ) );
  NOR2_X1 U1060 ( .A1(n116), .A2(n98), .ZN(\ab[4][11] ) );
  NOR2_X1 U1061 ( .A1(n190), .A2(n102), .ZN(\ab[6][9] ) );
  NOR2_X1 U1062 ( .A1(n184), .A2(n108), .ZN(\ab[8][7] ) );
  NOR2_X1 U1063 ( .A1(n180), .A2(n89), .ZN(\ab[10][5] ) );
  NOR2_X1 U1064 ( .A1(n172), .A2(n61), .ZN(\ab[15][2] ) );
  NOR2_X1 U1065 ( .A1(n116), .A2(n96), .ZN(\ab[3][11] ) );
  NOR2_X1 U1066 ( .A1(n116), .A2(net144909), .ZN(\ab[2][11] ) );
  AND2_X1 U1067 ( .A1(\ab[1][11] ), .A2(\ab[0][12] ), .ZN(\CARRYB[1][11] ) );
  NOR2_X1 U1068 ( .A1(n190), .A2(n99), .ZN(\ab[5][9] ) );
  NOR2_X1 U1069 ( .A1(n190), .A2(n97), .ZN(\ab[4][9] ) );
  NOR2_X1 U1070 ( .A1(n184), .A2(n105), .ZN(\ab[7][7] ) );
  NOR2_X1 U1071 ( .A1(n184), .A2(n102), .ZN(\ab[6][7] ) );
  NOR2_X1 U1072 ( .A1(n193), .A2(n178), .ZN(\ab[9][5] ) );
  NOR2_X1 U1073 ( .A1(n178), .A2(n108), .ZN(\ab[8][5] ) );
  NOR2_X1 U1074 ( .A1(n175), .A2(n93), .ZN(\ab[12][3] ) );
  NOR2_X1 U1075 ( .A1(n172), .A2(n62), .ZN(\ab[14][2] ) );
  NOR2_X1 U1076 ( .A1(n144), .A2(n57), .ZN(\ab[19][1] ) );
  NOR2_X1 U1077 ( .A1(n175), .A2(n65), .ZN(\ab[11][3] ) );
  NOR2_X1 U1078 ( .A1(n175), .A2(n89), .ZN(\ab[10][3] ) );
  NOR2_X1 U1079 ( .A1(n190), .A2(n95), .ZN(\ab[3][9] ) );
  NOR2_X1 U1080 ( .A1(n184), .A2(n99), .ZN(\ab[5][7] ) );
  NOR2_X1 U1081 ( .A1(n178), .A2(n105), .ZN(\ab[7][5] ) );
  NOR2_X1 U1082 ( .A1(n144), .A2(n58), .ZN(\ab[18][1] ) );
  NOR2_X1 U1083 ( .A1(n172), .A2(n63), .ZN(\ab[13][2] ) );
  NOR2_X1 U1084 ( .A1(n193), .A2(n173), .ZN(\ab[9][3] ) );
  NOR2_X1 U1085 ( .A1(n190), .A2(net144909), .ZN(\ab[2][9] ) );
  AND2_X1 U1086 ( .A1(\ab[1][9] ), .A2(\ab[0][10] ), .ZN(\CARRYB[1][9] ) );
  NOR2_X1 U1087 ( .A1(n184), .A2(n97), .ZN(\ab[4][7] ) );
  NOR2_X1 U1088 ( .A1(n178), .A2(n102), .ZN(\ab[6][5] ) );
  NOR2_X1 U1089 ( .A1(n144), .A2(n59), .ZN(\ab[17][1] ) );
  NOR2_X1 U1090 ( .A1(n172), .A2(n93), .ZN(\ab[12][2] ) );
  NOR2_X1 U1091 ( .A1(n172), .A2(n65), .ZN(\ab[11][2] ) );
  NOR2_X1 U1092 ( .A1(n145), .A2(n60), .ZN(\ab[16][1] ) );
  NOR2_X1 U1093 ( .A1(n173), .A2(n108), .ZN(\ab[8][3] ) );
  NOR2_X1 U1094 ( .A1(n172), .A2(n89), .ZN(\ab[10][2] ) );
  NOR2_X1 U1095 ( .A1(n145), .A2(n61), .ZN(\ab[15][1] ) );
  NOR2_X1 U1096 ( .A1(n184), .A2(n95), .ZN(\ab[3][7] ) );
  NOR2_X1 U1097 ( .A1(n184), .A2(net144909), .ZN(\ab[2][7] ) );
  AND2_X1 U1098 ( .A1(\ab[1][7] ), .A2(\ab[0][8] ), .ZN(\CARRYB[1][7] ) );
  NOR2_X1 U1099 ( .A1(n178), .A2(n99), .ZN(\ab[5][5] ) );
  NOR2_X1 U1100 ( .A1(n178), .A2(n97), .ZN(\ab[4][5] ) );
  NOR2_X1 U1101 ( .A1(n193), .A2(n171), .ZN(\ab[9][2] ) );
  NOR2_X1 U1102 ( .A1(n178), .A2(n96), .ZN(\ab[3][5] ) );
  NOR2_X1 U1103 ( .A1(n173), .A2(n105), .ZN(\ab[7][3] ) );
  NOR2_X1 U1104 ( .A1(n145), .A2(n62), .ZN(\ab[14][1] ) );
  NOR2_X1 U1105 ( .A1(n173), .A2(n102), .ZN(\ab[6][3] ) );
  NOR2_X1 U1106 ( .A1(n178), .A2(net144909), .ZN(\ab[2][5] ) );
  AND2_X1 U1107 ( .A1(\ab[1][5] ), .A2(\ab[0][6] ), .ZN(\CARRYB[1][5] ) );
  NOR2_X1 U1108 ( .A1(n145), .A2(n63), .ZN(\ab[13][1] ) );
  NOR2_X1 U1109 ( .A1(n173), .A2(n99), .ZN(\ab[5][3] ) );
  NOR2_X1 U1110 ( .A1(n145), .A2(n64), .ZN(\ab[12][1] ) );
  NOR2_X1 U1111 ( .A1(n171), .A2(n108), .ZN(\ab[8][2] ) );
  NOR2_X1 U1112 ( .A1(n173), .A2(n97), .ZN(\ab[4][3] ) );
  NOR2_X1 U1113 ( .A1(n145), .A2(n92), .ZN(\ab[11][1] ) );
  NOR2_X1 U1114 ( .A1(n171), .A2(n105), .ZN(\ab[7][2] ) );
  NOR2_X1 U1115 ( .A1(n171), .A2(n102), .ZN(\ab[6][2] ) );
  NOR2_X1 U1116 ( .A1(n173), .A2(n96), .ZN(\ab[3][3] ) );
  NOR2_X1 U1117 ( .A1(n145), .A2(n90), .ZN(\ab[10][1] ) );
  NOR2_X1 U1118 ( .A1(n171), .A2(n99), .ZN(\ab[5][2] ) );
  NOR2_X1 U1119 ( .A1(n173), .A2(net144909), .ZN(\ab[2][3] ) );
  AND2_X1 U1120 ( .A1(\ab[1][3] ), .A2(\ab[0][4] ), .ZN(\CARRYB[1][3] ) );
  NOR2_X1 U1121 ( .A1(n171), .A2(n97), .ZN(\ab[4][2] ) );
  NOR2_X1 U1122 ( .A1(n194), .A2(n143), .ZN(\ab[9][1] ) );
  NOR2_X1 U1123 ( .A1(n143), .A2(n109), .ZN(\ab[8][1] ) );
  NOR2_X1 U1124 ( .A1(n171), .A2(n95), .ZN(\ab[3][2] ) );
  NOR2_X1 U1125 ( .A1(n143), .A2(n106), .ZN(\ab[7][1] ) );
  NOR2_X1 U1126 ( .A1(n171), .A2(n45), .ZN(\ab[2][2] ) );
  AND2_X1 U1127 ( .A1(\ab[1][2] ), .A2(\ab[0][3] ), .ZN(\CARRYB[1][2] ) );
  NOR2_X1 U1128 ( .A1(n143), .A2(n103), .ZN(\ab[6][1] ) );
  NOR2_X1 U1129 ( .A1(n143), .A2(n100), .ZN(\ab[5][1] ) );
  NOR2_X1 U1130 ( .A1(n143), .A2(n98), .ZN(\ab[4][1] ) );
  NOR2_X1 U1131 ( .A1(n143), .A2(n96), .ZN(\ab[3][1] ) );
  NOR2_X1 U1132 ( .A1(n143), .A2(net144909), .ZN(\ab[2][1] ) );
  AND2_X1 U1133 ( .A1(\ab[1][1] ), .A2(\ab[0][2] ), .ZN(\CARRYB[1][1] ) );
  NOR2_X1 U1134 ( .A1(n111), .A2(n46), .ZN(\ab[29][0] ) );
  NOR2_X1 U1135 ( .A1(n111), .A2(n44), .ZN(\ab[30][0] ) );
  NOR2_X1 U1136 ( .A1(n111), .A2(n47), .ZN(\ab[28][0] ) );
  NOR2_X1 U1137 ( .A1(n112), .A2(n48), .ZN(\ab[27][0] ) );
  NOR2_X1 U1138 ( .A1(n112), .A2(n49), .ZN(\ab[26][0] ) );
  NOR2_X1 U1139 ( .A1(n112), .A2(n50), .ZN(\ab[25][0] ) );
  NOR2_X1 U1140 ( .A1(n112), .A2(n51), .ZN(\ab[24][0] ) );
  NOR2_X1 U1141 ( .A1(n112), .A2(n52), .ZN(\ab[23][0] ) );
  NOR2_X1 U1142 ( .A1(n112), .A2(n53), .ZN(\ab[22][0] ) );
  NOR2_X1 U1143 ( .A1(n112), .A2(n54), .ZN(\ab[21][0] ) );
  NOR2_X1 U1144 ( .A1(n112), .A2(n55), .ZN(\ab[20][0] ) );
  NOR2_X1 U1145 ( .A1(n112), .A2(n57), .ZN(\ab[19][0] ) );
  NOR2_X1 U1146 ( .A1(n112), .A2(n58), .ZN(\ab[18][0] ) );
  NOR2_X1 U1147 ( .A1(n112), .A2(n59), .ZN(\ab[17][0] ) );
  NOR2_X1 U1148 ( .A1(n112), .A2(n60), .ZN(\ab[16][0] ) );
  NOR2_X1 U1149 ( .A1(n112), .A2(n61), .ZN(\ab[15][0] ) );
  NOR2_X1 U1150 ( .A1(n112), .A2(n62), .ZN(\ab[14][0] ) );
  NOR2_X1 U1151 ( .A1(n112), .A2(n63), .ZN(\ab[13][0] ) );
  NOR2_X1 U1152 ( .A1(n112), .A2(n64), .ZN(\ab[12][0] ) );
  NOR2_X1 U1153 ( .A1(n112), .A2(n65), .ZN(\ab[11][0] ) );
  NOR2_X1 U1154 ( .A1(n172), .A2(net145039), .ZN(\ab[0][2] ) );
  NOR2_X1 U1155 ( .A1(n145), .A2(net145041), .ZN(\ab[0][1] ) );
  NOR2_X1 U1156 ( .A1(n36), .A2(net144973), .ZN(\ab[1][0] ) );
  NOR2_X1 U1157 ( .A1(net144707), .A2(n44), .ZN(\ab[30][31] ) );
  NOR2_X1 U1158 ( .A1(net144717), .A2(n43), .ZN(\ab[31][30] ) );
  NOR2_X1 U1159 ( .A1(n170), .A2(n43), .ZN(\ab[31][29] ) );
  NOR2_X1 U1160 ( .A1(n161), .A2(n43), .ZN(\ab[31][25] ) );
  NOR2_X1 U1161 ( .A1(n160), .A2(n43), .ZN(\ab[31][24] ) );
  NOR2_X1 U1162 ( .A1(n164), .A2(n43), .ZN(\ab[31][26] ) );
  NOR2_X1 U1163 ( .A1(n157), .A2(n43), .ZN(\ab[31][23] ) );
  NOR2_X1 U1164 ( .A1(n166), .A2(n43), .ZN(\ab[31][27] ) );
  NOR2_X1 U1165 ( .A1(n152), .A2(n43), .ZN(\ab[31][22] ) );
  NOR2_X1 U1166 ( .A1(n151), .A2(n43), .ZN(\ab[31][21] ) );
  NOR2_X1 U1167 ( .A1(n168), .A2(n43), .ZN(\ab[31][28] ) );
  NOR2_X1 U1168 ( .A1(n146), .A2(n43), .ZN(\ab[31][20] ) );
  NOR2_X1 U1169 ( .A1(n140), .A2(n43), .ZN(\ab[31][19] ) );
  NOR2_X1 U1170 ( .A1(n137), .A2(n43), .ZN(\ab[31][18] ) );
  NOR2_X1 U1171 ( .A1(n134), .A2(n43), .ZN(\ab[31][17] ) );
  NOR2_X1 U1172 ( .A1(n144), .A2(n79), .ZN(\ab[1][1] ) );
  NOR2_X1 U1173 ( .A1(net169601), .A2(n44), .ZN(\ab[30][30] ) );
  NOR2_X1 U1174 ( .A1(net144709), .A2(n46), .ZN(\ab[29][31] ) );
  NOR2_X1 U1175 ( .A1(net144709), .A2(n59), .ZN(\ab[17][31] ) );
  NOR2_X1 U1176 ( .A1(net169601), .A2(n58), .ZN(\ab[18][30] ) );
  NOR2_X1 U1177 ( .A1(net144707), .A2(n58), .ZN(\ab[18][31] ) );
  NOR2_X1 U1178 ( .A1(net144717), .A2(n57), .ZN(\ab[19][30] ) );
  NOR2_X1 U1179 ( .A1(net144709), .A2(n57), .ZN(\ab[19][31] ) );
  NOR2_X1 U1180 ( .A1(net169601), .A2(n55), .ZN(\ab[20][30] ) );
  NOR2_X1 U1181 ( .A1(net144707), .A2(n55), .ZN(\ab[20][31] ) );
  NOR2_X1 U1182 ( .A1(net144717), .A2(n54), .ZN(\ab[21][30] ) );
  NOR2_X1 U1183 ( .A1(net144709), .A2(n54), .ZN(\ab[21][31] ) );
  NOR2_X1 U1184 ( .A1(net169601), .A2(n53), .ZN(\ab[22][30] ) );
  NOR2_X1 U1185 ( .A1(net144707), .A2(n53), .ZN(\ab[22][31] ) );
  NOR2_X1 U1186 ( .A1(net144717), .A2(n52), .ZN(\ab[23][30] ) );
  NOR2_X1 U1187 ( .A1(net169601), .A2(n51), .ZN(\ab[24][30] ) );
  NOR2_X1 U1188 ( .A1(net144709), .A2(n52), .ZN(\ab[23][31] ) );
  NOR2_X1 U1189 ( .A1(net144707), .A2(n51), .ZN(\ab[24][31] ) );
  NOR2_X1 U1190 ( .A1(net144717), .A2(n50), .ZN(\ab[25][30] ) );
  NOR2_X1 U1191 ( .A1(net169601), .A2(n49), .ZN(\ab[26][30] ) );
  NOR2_X1 U1192 ( .A1(net144709), .A2(n50), .ZN(\ab[25][31] ) );
  NOR2_X1 U1193 ( .A1(net144707), .A2(n49), .ZN(\ab[26][31] ) );
  NOR2_X1 U1194 ( .A1(net144717), .A2(n48), .ZN(\ab[27][30] ) );
  NOR2_X1 U1195 ( .A1(net144717), .A2(n46), .ZN(\ab[29][30] ) );
  NOR2_X1 U1196 ( .A1(net144707), .A2(n47), .ZN(\ab[28][31] ) );
  NOR2_X1 U1197 ( .A1(net144709), .A2(n48), .ZN(\ab[27][31] ) );
  NOR2_X1 U1198 ( .A1(net169601), .A2(n47), .ZN(\ab[28][30] ) );
  NOR2_X1 U1199 ( .A1(n162), .A2(n44), .ZN(\ab[30][25] ) );
  NOR2_X1 U1200 ( .A1(n158), .A2(n44), .ZN(\ab[30][24] ) );
  NOR2_X1 U1201 ( .A1(n155), .A2(n44), .ZN(\ab[30][23] ) );
  NOR2_X1 U1202 ( .A1(n163), .A2(n44), .ZN(\ab[30][26] ) );
  NOR2_X1 U1203 ( .A1(n152), .A2(n44), .ZN(\ab[30][22] ) );
  NOR2_X1 U1204 ( .A1(n167), .A2(n44), .ZN(\ab[30][27] ) );
  NOR2_X1 U1205 ( .A1(n150), .A2(n44), .ZN(\ab[30][21] ) );
  NOR2_X1 U1206 ( .A1(n160), .A2(n46), .ZN(\ab[29][24] ) );
  NOR2_X1 U1207 ( .A1(n162), .A2(n46), .ZN(\ab[29][25] ) );
  NOR2_X1 U1208 ( .A1(n146), .A2(n44), .ZN(\ab[30][20] ) );
  NOR2_X1 U1209 ( .A1(n157), .A2(n46), .ZN(\ab[29][23] ) );
  NOR2_X1 U1210 ( .A1(n164), .A2(n46), .ZN(\ab[29][26] ) );
  NOR2_X1 U1211 ( .A1(n152), .A2(n46), .ZN(\ab[29][22] ) );
  NOR2_X1 U1212 ( .A1(n140), .A2(n44), .ZN(\ab[30][19] ) );
  NOR2_X1 U1213 ( .A1(n168), .A2(n44), .ZN(\ab[30][28] ) );
  NOR2_X1 U1214 ( .A1(n149), .A2(n46), .ZN(\ab[29][21] ) );
  NOR2_X1 U1215 ( .A1(n166), .A2(n46), .ZN(\ab[29][27] ) );
  NOR2_X1 U1218 ( .A1(n137), .A2(n44), .ZN(\ab[30][18] ) );
  NOR2_X1 U1219 ( .A1(n146), .A2(n46), .ZN(\ab[29][20] ) );
  NOR2_X1 U1220 ( .A1(n158), .A2(n47), .ZN(\ab[28][24] ) );
  NOR2_X1 U1221 ( .A1(n161), .A2(n47), .ZN(\ab[28][25] ) );
  NOR2_X1 U1222 ( .A1(n170), .A2(n44), .ZN(\ab[30][29] ) );
  NOR2_X1 U1223 ( .A1(n155), .A2(n47), .ZN(\ab[28][23] ) );
  NOR2_X1 U1224 ( .A1(n140), .A2(n46), .ZN(\ab[29][19] ) );
  NOR2_X1 U1225 ( .A1(n152), .A2(n47), .ZN(\ab[28][22] ) );
  NOR2_X1 U1226 ( .A1(n163), .A2(n47), .ZN(\ab[28][26] ) );
  NOR2_X1 U1227 ( .A1(n151), .A2(n47), .ZN(\ab[28][21] ) );
  NOR2_X1 U1228 ( .A1(n146), .A2(n47), .ZN(\ab[28][20] ) );
  NOR2_X1 U1229 ( .A1(n153), .A2(n49), .ZN(\ab[26][22] ) );
  NOR2_X1 U1230 ( .A1(n158), .A2(n51), .ZN(\ab[24][24] ) );
  NOR2_X1 U1231 ( .A1(n163), .A2(n53), .ZN(\ab[22][26] ) );
  NOR2_X1 U1232 ( .A1(n169), .A2(n55), .ZN(\ab[20][28] ) );
  NOR2_X1 U1233 ( .A1(n150), .A2(n48), .ZN(\ab[27][21] ) );
  NOR2_X1 U1234 ( .A1(n157), .A2(n50), .ZN(\ab[25][23] ) );
  NOR2_X1 U1235 ( .A1(n162), .A2(n52), .ZN(\ab[23][25] ) );
  NOR2_X1 U1236 ( .A1(n166), .A2(n54), .ZN(\ab[21][27] ) );
  NOR2_X1 U1237 ( .A1(n170), .A2(n57), .ZN(\ab[19][29] ) );
  NOR2_X1 U1238 ( .A1(n169), .A2(n46), .ZN(\ab[29][28] ) );
  NOR2_X1 U1239 ( .A1(n155), .A2(n49), .ZN(\ab[26][23] ) );
  NOR2_X1 U1240 ( .A1(n162), .A2(n51), .ZN(\ab[24][25] ) );
  NOR2_X1 U1241 ( .A1(n167), .A2(n53), .ZN(\ab[22][27] ) );
  NOR2_X1 U1242 ( .A1(n170), .A2(n55), .ZN(\ab[20][29] ) );
  NOR2_X1 U1243 ( .A1(n153), .A2(n48), .ZN(\ab[27][22] ) );
  NOR2_X1 U1244 ( .A1(n158), .A2(n50), .ZN(\ab[25][24] ) );
  NOR2_X1 U1245 ( .A1(n164), .A2(n52), .ZN(\ab[23][26] ) );
  NOR2_X1 U1246 ( .A1(n168), .A2(n54), .ZN(\ab[21][28] ) );
  NOR2_X1 U1247 ( .A1(n167), .A2(n47), .ZN(\ab[28][27] ) );
  NOR2_X1 U1248 ( .A1(n157), .A2(n48), .ZN(\ab[27][23] ) );
  NOR2_X1 U1249 ( .A1(n161), .A2(n50), .ZN(\ab[25][25] ) );
  NOR2_X1 U1250 ( .A1(n166), .A2(n52), .ZN(\ab[23][27] ) );
  NOR2_X1 U1251 ( .A1(n170), .A2(n54), .ZN(\ab[21][29] ) );
  NOR2_X1 U1252 ( .A1(n160), .A2(n49), .ZN(\ab[26][24] ) );
  NOR2_X1 U1253 ( .A1(n163), .A2(n51), .ZN(\ab[24][26] ) );
  NOR2_X1 U1254 ( .A1(n169), .A2(n53), .ZN(\ab[22][28] ) );
  NOR2_X1 U1255 ( .A1(n158), .A2(n48), .ZN(\ab[27][24] ) );
  NOR2_X1 U1256 ( .A1(n162), .A2(n49), .ZN(\ab[26][25] ) );
  NOR2_X1 U1257 ( .A1(n167), .A2(n51), .ZN(\ab[24][27] ) );
  NOR2_X1 U1258 ( .A1(n170), .A2(n53), .ZN(\ab[22][29] ) );
  NOR2_X1 U1259 ( .A1(n163), .A2(n50), .ZN(\ab[25][26] ) );
  NOR2_X1 U1260 ( .A1(n169), .A2(n52), .ZN(\ab[23][28] ) );
  NOR2_X1 U1261 ( .A1(n162), .A2(n48), .ZN(\ab[27][25] ) );
  NOR2_X1 U1262 ( .A1(n166), .A2(n50), .ZN(\ab[25][27] ) );
  NOR2_X1 U1263 ( .A1(n170), .A2(n52), .ZN(\ab[23][29] ) );
  NOR2_X1 U1264 ( .A1(n164), .A2(n49), .ZN(\ab[26][26] ) );
  NOR2_X1 U1265 ( .A1(n168), .A2(n51), .ZN(\ab[24][28] ) );
  NOR2_X1 U1266 ( .A1(n163), .A2(n48), .ZN(\ab[27][26] ) );
  NOR2_X1 U1267 ( .A1(n167), .A2(n49), .ZN(\ab[26][27] ) );
  NOR2_X1 U1268 ( .A1(n170), .A2(n51), .ZN(\ab[24][29] ) );
  NOR2_X1 U1269 ( .A1(n169), .A2(n50), .ZN(\ab[25][28] ) );
  NOR2_X1 U1270 ( .A1(n166), .A2(n48), .ZN(\ab[27][27] ) );
  NOR2_X1 U1271 ( .A1(n170), .A2(n50), .ZN(\ab[25][29] ) );
  NOR2_X1 U1272 ( .A1(n168), .A2(n49), .ZN(\ab[26][28] ) );
  NOR2_X1 U1273 ( .A1(n168), .A2(n47), .ZN(\ab[28][28] ) );
  NOR2_X1 U1274 ( .A1(n169), .A2(n48), .ZN(\ab[27][28] ) );
  NOR2_X1 U1275 ( .A1(n170), .A2(n49), .ZN(\ab[26][29] ) );
  NOR2_X1 U1276 ( .A1(n170), .A2(n46), .ZN(\ab[29][29] ) );
  NOR2_X1 U1277 ( .A1(n170), .A2(n48), .ZN(\ab[27][29] ) );
  NOR2_X1 U1278 ( .A1(n170), .A2(n47), .ZN(\ab[28][29] ) );
  NOR2_X1 U1279 ( .A1(n112), .A2(n91), .ZN(\ab[10][0] ) );
  NOR2_X1 U1280 ( .A1(n195), .A2(n111), .ZN(\ab[9][0] ) );
  NOR2_X1 U1281 ( .A1(n111), .A2(n110), .ZN(\ab[8][0] ) );
  NOR2_X1 U1282 ( .A1(n111), .A2(n107), .ZN(\ab[7][0] ) );
  NOR2_X1 U1283 ( .A1(n111), .A2(n104), .ZN(\ab[6][0] ) );
  NOR2_X1 U1284 ( .A1(n111), .A2(n101), .ZN(\ab[5][0] ) );
  NOR2_X1 U1285 ( .A1(n111), .A2(n41), .ZN(\ab[4][0] ) );
  NOR2_X1 U1286 ( .A1(n111), .A2(n45), .ZN(\ab[2][0] ) );
  AND2_X1 U1287 ( .A1(\ab[1][0] ), .A2(\ab[0][1] ), .ZN(\CARRYB[1][0] ) );
  NOR2_X1 U1288 ( .A1(n111), .A2(n95), .ZN(\ab[3][0] ) );
  NOR2_X1 U1289 ( .A1(net144709), .A2(n43), .ZN(\SUMB[31][31] ) );
  NOR2_X1 U1290 ( .A1(n112), .A2(net145039), .ZN(PRODUCT[0]) );
  BUF_X2 U1291 ( .A(n23), .Z(n149) );
  BUF_X1 U1292 ( .A(n22), .Z(n154) );
  BUF_X1 U1293 ( .A(n24), .Z(n148) );
  BUF_X1 U1294 ( .A(n26), .Z(n142) );
  BUF_X1 U1295 ( .A(n27), .Z(n139) );
  BUF_X1 U1296 ( .A(n28), .Z(n136) );
  BUF_X1 U1297 ( .A(n29), .Z(n133) );
  BUF_X1 U1298 ( .A(n30), .Z(n130) );
  BUF_X1 U1299 ( .A(n32), .Z(n124) );
  BUF_X1 U1300 ( .A(n31), .Z(n127) );
  BUF_X1 U1301 ( .A(n33), .Z(n121) );
  BUF_X1 U1302 ( .A(n34), .Z(n118) );
  BUF_X1 U1303 ( .A(n35), .Z(n115) );
  BUF_X1 U1304 ( .A(n5), .Z(n192) );
  BUF_X1 U1305 ( .A(n6), .Z(n189) );
  BUF_X1 U1306 ( .A(n7), .Z(n186) );
  BUF_X1 U1307 ( .A(n8), .Z(n183) );
  BUF_X1 U1308 ( .A(n9), .Z(n180) );
  BUF_X1 U1309 ( .A(n10), .Z(n177) );
  BUF_X1 U1310 ( .A(n11), .Z(n175) );
  BUF_X1 U1311 ( .A(n66), .Z(n90) );
  BUF_X1 U1312 ( .A(n66), .Z(n89) );
  BUF_X1 U1313 ( .A(n40), .Z(n101) );
  BUF_X1 U1314 ( .A(n39), .Z(n104) );
  BUF_X1 U1315 ( .A(n38), .Z(n107) );
  BUF_X1 U1316 ( .A(n37), .Z(n110) );
  BUF_X1 U1317 ( .A(n25), .Z(n145) );
  BUF_X1 U1318 ( .A(n4), .Z(n195) );
  CLKBUF_X1 U1319 ( .A(n36), .Z(n112) );
  INV_X1 U1320 ( .A(B[25]), .ZN(n19) );
  INV_X1 U1321 ( .A(B[26]), .ZN(n18) );
  INV_X1 U1322 ( .A(B[24]), .ZN(n20) );
  INV_X1 U1323 ( .A(B[27]), .ZN(n17) );
  INV_X1 U1324 ( .A(B[23]), .ZN(n21) );
  INV_X1 U1325 ( .A(B[22]), .ZN(n22) );
  INV_X1 U1326 ( .A(B[28]), .ZN(n16) );
  INV_X1 U1327 ( .A(B[21]), .ZN(n23) );
  INV_X1 U1328 ( .A(B[20]), .ZN(n24) );
  INV_X1 U1329 ( .A(B[19]), .ZN(n26) );
  INV_X1 U1330 ( .A(B[18]), .ZN(n27) );
  INV_X1 U1331 ( .A(B[17]), .ZN(n28) );
  INV_X1 U1332 ( .A(B[16]), .ZN(n29) );
  INV_X1 U1333 ( .A(B[15]), .ZN(n30) );
  INV_X1 U1334 ( .A(B[12]), .ZN(n33) );
  INV_X1 U1335 ( .A(B[13]), .ZN(n32) );
  INV_X1 U1336 ( .A(B[11]), .ZN(n34) );
  INV_X1 U1337 ( .A(B[14]), .ZN(n31) );
  INV_X1 U1338 ( .A(B[10]), .ZN(n35) );
  INV_X1 U1339 ( .A(A[3]), .ZN(n42) );
  INV_X1 U1340 ( .A(B[8]), .ZN(n6) );
  INV_X1 U1341 ( .A(B[7]), .ZN(n7) );
  INV_X1 U1342 ( .A(A[4]), .ZN(n41) );
  INV_X1 U1343 ( .A(B[6]), .ZN(n8) );
  INV_X1 U1344 ( .A(B[5]), .ZN(n9) );
  INV_X1 U1345 ( .A(B[3]), .ZN(n11) );
  INV_X1 U1346 ( .A(A[5]), .ZN(n40) );
  INV_X1 U1347 ( .A(A[6]), .ZN(n39) );
  INV_X1 U1348 ( .A(B[9]), .ZN(n5) );
  INV_X1 U1349 ( .A(B[1]), .ZN(n25) );
  INV_X1 U1350 ( .A(B[0]), .ZN(n36) );
  INV_X1 U1351 ( .A(A[10]), .ZN(n66) );
  INV_X1 U1352 ( .A(A[7]), .ZN(n38) );
  INV_X1 U1353 ( .A(A[8]), .ZN(n37) );
  INV_X1 U1354 ( .A(A[9]), .ZN(n4) );
  NOR2_X1 U1355 ( .A1(n14), .A2(net144973), .ZN(\ab[1][2] ) );
  NOR2_X1 U1356 ( .A1(n174), .A2(n79), .ZN(\ab[1][3] ) );
  NOR2_X1 U1357 ( .A1(n10), .A2(net144973), .ZN(\ab[1][4] ) );
  NOR2_X1 U1358 ( .A1(n179), .A2(net144973), .ZN(\ab[1][5] ) );
  NOR2_X1 U1359 ( .A1(n182), .A2(n79), .ZN(\ab[1][6] ) );
  NOR2_X1 U1360 ( .A1(n185), .A2(net144973), .ZN(\ab[1][7] ) );
  NOR2_X1 U1361 ( .A1(n188), .A2(n79), .ZN(\ab[1][8] ) );
  NOR2_X1 U1362 ( .A1(n191), .A2(net144973), .ZN(\ab[1][9] ) );
  NOR2_X1 U1363 ( .A1(n56), .A2(n15), .ZN(\ab[1][29] ) );
endmodule


module Flag_Generator_NBIT_ALU32 ( FG_ALU_out, FG_sgn_usgn, FG_carry, FG_ZF, 
        FG_PF, FG_SF, FG_CF, FG_OF );
  input [31:0] FG_ALU_out;
  input FG_sgn_usgn, FG_carry;
  output FG_ZF, FG_PF, FG_SF, FG_CF, FG_OF;
  wire   n2, n3;

  NORGate_NX1_N32 NOR32X1 ( .A({FG_ALU_out[31:1], n3}), .B({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y(FG_ZF) );
  XNORGate_NX1_N32 XNOR32X1 ( .A(FG_ALU_out), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .Y(FG_PF) );
  CLKBUF_X1 U2 ( .A(FG_ALU_out[0]), .Z(n3) );
  NOR2_X1 U3 ( .A1(FG_sgn_usgn), .A2(n2), .ZN(FG_CF) );
  INV_X1 U4 ( .A(FG_carry), .ZN(n2) );
  AND2_X1 U5 ( .A1(FG_sgn_usgn), .A2(FG_ALU_out[31]), .ZN(FG_SF) );
  AND2_X1 U6 ( .A1(FG_sgn_usgn), .A2(FG_carry), .ZN(FG_OF) );
endmodule


module Comparison_Logic_NBIT_DATA32 ( CMPL_OpA, CMPL_OpB, CMPL_OPCODE, CMPL_Y
 );
  input [31:0] CMPL_OpA;
  input [31:0] CMPL_OpB;
  input [3:0] CMPL_OPCODE;
  output [31:0] CMPL_Y;
  wire   s_A_gt_B, s_A_ge_B, s_A_lt_B, s_A_le_B, s_A_eq_B, n4, n5, n6, n7, n8,
         n9, n10, n11, n12;
  assign CMPL_Y[31] = 1'b0;
  assign CMPL_Y[30] = 1'b0;
  assign CMPL_Y[29] = 1'b0;
  assign CMPL_Y[28] = 1'b0;
  assign CMPL_Y[27] = 1'b0;
  assign CMPL_Y[26] = 1'b0;
  assign CMPL_Y[25] = 1'b0;
  assign CMPL_Y[24] = 1'b0;
  assign CMPL_Y[23] = 1'b0;
  assign CMPL_Y[22] = 1'b0;
  assign CMPL_Y[21] = 1'b0;
  assign CMPL_Y[20] = 1'b0;
  assign CMPL_Y[19] = 1'b0;
  assign CMPL_Y[18] = 1'b0;
  assign CMPL_Y[17] = 1'b0;
  assign CMPL_Y[16] = 1'b0;
  assign CMPL_Y[15] = 1'b0;
  assign CMPL_Y[14] = 1'b0;
  assign CMPL_Y[13] = 1'b0;
  assign CMPL_Y[12] = 1'b0;
  assign CMPL_Y[11] = 1'b0;
  assign CMPL_Y[10] = 1'b0;
  assign CMPL_Y[9] = 1'b0;
  assign CMPL_Y[8] = 1'b0;
  assign CMPL_Y[7] = 1'b0;
  assign CMPL_Y[6] = 1'b0;
  assign CMPL_Y[5] = 1'b0;
  assign CMPL_Y[4] = 1'b0;
  assign CMPL_Y[3] = 1'b0;
  assign CMPL_Y[2] = 1'b0;
  assign CMPL_Y[1] = 1'b0;

  NAND3_X1 U10 ( .A1(n6), .A2(n7), .A3(CMPL_OPCODE[2]), .ZN(n5) );
  XOR2_X1 U11 ( .A(s_A_eq_B), .B(CMPL_OPCODE[0]), .Z(n6) );
  Comparator_NBIT_DATA32 CMP ( .CMP_OpA(CMPL_OpA), .CMP_OpB(CMPL_OpB), 
        .CMP_sgn_usgn(CMPL_OPCODE[3]), .CMP_A_gt_B(s_A_gt_B), .CMP_A_ge_B(
        s_A_ge_B), .CMP_A_lt_B(s_A_lt_B), .CMP_A_le_B(s_A_le_B), .CMP_A_eq_B(
        s_A_eq_B) );
  INV_X1 U2 ( .A(CMPL_OPCODE[1]), .ZN(n7) );
  INV_X1 U3 ( .A(CMPL_OPCODE[0]), .ZN(n12) );
  INV_X1 U4 ( .A(CMPL_OPCODE[2]), .ZN(n9) );
  AOI22_X1 U5 ( .A1(s_A_lt_B), .A2(n12), .B1(s_A_gt_B), .B2(CMPL_OPCODE[0]), 
        .ZN(n11) );
  NAND2_X1 U6 ( .A1(n4), .A2(n5), .ZN(CMPL_Y[0]) );
  OAI22_X1 U7 ( .A1(n10), .A2(n7), .B1(CMPL_OPCODE[1]), .B2(n11), .ZN(n8) );
  AOI22_X1 U8 ( .A1(s_A_le_B), .A2(n12), .B1(s_A_ge_B), .B2(CMPL_OPCODE[0]), 
        .ZN(n10) );
  NAND2_X1 U9 ( .A1(n8), .A2(n9), .ZN(n4) );
endmodule


module Logic_Unit_NBIT_DATA32 ( LU_OpA, LU_OpB, LU_Opcode, LU_Y );
  input [31:0] LU_OpA;
  input [31:0] LU_OpB;
  input [3:0] LU_Opcode;
  output [31:0] LU_Y;
  wire   n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78,
         n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92,
         n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, n135, n136, n137, n138,
         n139, n140, n141, n142, n143, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n175, n176, n177, n178, n179, n180, n181, n182,
         n183, n184, n185, n186, n187, n188, n189, n190, n191, n192, n193,
         n194, n195, n196, n197, n198, n199, n200, n201, n202, n203, n204;

  INV_X1 U1 ( .A(LU_OpA[21]), .ZN(n140) );
  INV_X1 U2 ( .A(LU_OpA[18]), .ZN(n156) );
  INV_X1 U3 ( .A(LU_OpA[3]), .ZN(n92) );
  INV_X1 U4 ( .A(LU_OpA[24]), .ZN(n128) );
  INV_X1 U5 ( .A(LU_OpA[27]), .ZN(n116) );
  INV_X1 U6 ( .A(LU_OpA[9]), .ZN(n68) );
  INV_X1 U7 ( .A(LU_OpA[12]), .ZN(n180) );
  INV_X1 U8 ( .A(LU_OpA[15]), .ZN(n168) );
  INV_X1 U9 ( .A(LU_OpA[6]), .ZN(n80) );
  INV_X1 U10 ( .A(LU_OpA[1]), .ZN(n148) );
  INV_X1 U11 ( .A(LU_OpA[5]), .ZN(n84) );
  INV_X1 U12 ( .A(LU_OpA[16]), .ZN(n164) );
  INV_X1 U13 ( .A(LU_OpA[0]), .ZN(n192) );
  INV_X1 U14 ( .A(LU_OpA[11]), .ZN(n184) );
  INV_X1 U15 ( .A(LU_OpA[20]), .ZN(n144) );
  INV_X1 U16 ( .A(LU_OpA[23]), .ZN(n132) );
  INV_X1 U17 ( .A(LU_OpA[17]), .ZN(n160) );
  INV_X1 U18 ( .A(LU_OpA[14]), .ZN(n172) );
  INV_X1 U19 ( .A(LU_OpA[26]), .ZN(n120) );
  INV_X1 U20 ( .A(LU_OpA[8]), .ZN(n72) );
  INV_X1 U21 ( .A(LU_OpA[7]), .ZN(n76) );
  INV_X1 U22 ( .A(LU_OpA[4]), .ZN(n88) );
  INV_X1 U23 ( .A(LU_OpA[2]), .ZN(n104) );
  INV_X1 U24 ( .A(LU_OpA[28]), .ZN(n112) );
  INV_X1 U25 ( .A(LU_OpA[10]), .ZN(n188) );
  INV_X1 U26 ( .A(LU_OpA[19]), .ZN(n152) );
  INV_X1 U27 ( .A(LU_OpA[13]), .ZN(n176) );
  INV_X1 U28 ( .A(LU_OpA[29]), .ZN(n108) );
  INV_X1 U29 ( .A(LU_OpA[22]), .ZN(n136) );
  INV_X1 U30 ( .A(LU_OpA[25]), .ZN(n124) );
  OAI22_X1 U31 ( .A1(n97), .A2(n98), .B1(LU_OpB[30]), .B2(n99), .ZN(LU_Y[30])
         );
  INV_X1 U32 ( .A(LU_OpB[30]), .ZN(n98) );
  OAI22_X1 U33 ( .A1(n73), .A2(n74), .B1(LU_OpB[7]), .B2(n75), .ZN(LU_Y[7]) );
  INV_X1 U34 ( .A(LU_OpB[7]), .ZN(n74) );
  OAI22_X1 U35 ( .A1(n93), .A2(n94), .B1(LU_OpB[31]), .B2(n95), .ZN(LU_Y[31])
         );
  INV_X1 U36 ( .A(LU_OpB[31]), .ZN(n94) );
  OAI22_X1 U37 ( .A1(n185), .A2(n186), .B1(LU_OpB[10]), .B2(n187), .ZN(
        LU_Y[10]) );
  INV_X1 U38 ( .A(LU_OpB[10]), .ZN(n186) );
  OAI22_X1 U39 ( .A1(n181), .A2(n182), .B1(LU_OpB[11]), .B2(n183), .ZN(
        LU_Y[11]) );
  INV_X1 U40 ( .A(LU_OpB[11]), .ZN(n182) );
  OAI22_X1 U41 ( .A1(n133), .A2(n134), .B1(LU_OpB[22]), .B2(n135), .ZN(
        LU_Y[22]) );
  INV_X1 U42 ( .A(LU_OpB[22]), .ZN(n134) );
  OAI22_X1 U43 ( .A1(n129), .A2(n130), .B1(LU_OpB[23]), .B2(n131), .ZN(
        LU_Y[23]) );
  INV_X1 U44 ( .A(LU_OpB[23]), .ZN(n130) );
  OAI22_X1 U45 ( .A1(n153), .A2(n154), .B1(LU_OpB[18]), .B2(n155), .ZN(
        LU_Y[18]) );
  INV_X1 U46 ( .A(LU_OpB[18]), .ZN(n154) );
  OAI22_X1 U47 ( .A1(n149), .A2(n150), .B1(LU_OpB[19]), .B2(n151), .ZN(
        LU_Y[19]) );
  INV_X1 U48 ( .A(LU_OpB[19]), .ZN(n150) );
  OAI22_X1 U49 ( .A1(n169), .A2(n170), .B1(LU_OpB[14]), .B2(n171), .ZN(
        LU_Y[14]) );
  INV_X1 U50 ( .A(LU_OpB[14]), .ZN(n170) );
  OAI22_X1 U51 ( .A1(n165), .A2(n166), .B1(LU_OpB[15]), .B2(n167), .ZN(
        LU_Y[15]) );
  INV_X1 U52 ( .A(LU_OpB[15]), .ZN(n166) );
  OAI22_X1 U53 ( .A1(n117), .A2(n118), .B1(LU_OpB[26]), .B2(n119), .ZN(
        LU_Y[26]) );
  INV_X1 U54 ( .A(LU_OpB[26]), .ZN(n118) );
  OAI22_X1 U55 ( .A1(n113), .A2(n114), .B1(LU_OpB[27]), .B2(n115), .ZN(
        LU_Y[27]) );
  INV_X1 U56 ( .A(LU_OpB[27]), .ZN(n114) );
  OAI22_X1 U57 ( .A1(n89), .A2(n90), .B1(LU_OpB[3]), .B2(n91), .ZN(LU_Y[3]) );
  INV_X1 U58 ( .A(LU_OpB[3]), .ZN(n90) );
  OAI22_X1 U59 ( .A1(n77), .A2(n78), .B1(LU_OpB[6]), .B2(n79), .ZN(LU_Y[6]) );
  INV_X1 U60 ( .A(LU_OpB[6]), .ZN(n78) );
  AOI22_X1 U61 ( .A1(n195), .A2(n92), .B1(LU_OpA[3]), .B2(n201), .ZN(n91) );
  AOI22_X1 U62 ( .A1(n195), .A2(n88), .B1(LU_OpA[4]), .B2(n201), .ZN(n87) );
  AOI22_X1 U63 ( .A1(n195), .A2(n84), .B1(LU_OpA[5]), .B2(n201), .ZN(n83) );
  AOI22_X1 U64 ( .A1(n195), .A2(n72), .B1(LU_OpA[8]), .B2(n201), .ZN(n71) );
  AOI22_X1 U65 ( .A1(n195), .A2(n76), .B1(LU_OpA[7]), .B2(n201), .ZN(n75) );
  AOI22_X1 U66 ( .A1(n195), .A2(n80), .B1(LU_OpA[6]), .B2(n201), .ZN(n79) );
  AOI22_X1 U67 ( .A1(n195), .A2(n68), .B1(n201), .B2(LU_OpA[9]), .ZN(n67) );
  AOI22_X1 U68 ( .A1(n193), .A2(n192), .B1(LU_OpA[0]), .B2(n199), .ZN(n191) );
  AOI22_X1 U69 ( .A1(n193), .A2(n180), .B1(LU_OpA[12]), .B2(n199), .ZN(n179)
         );
  AOI22_X1 U70 ( .A1(n193), .A2(n188), .B1(LU_OpA[10]), .B2(n199), .ZN(n187)
         );
  AOI22_X1 U71 ( .A1(n193), .A2(n184), .B1(LU_OpA[11]), .B2(n199), .ZN(n183)
         );
  AOI22_X1 U72 ( .A1(n194), .A2(n144), .B1(LU_OpA[20]), .B2(n200), .ZN(n143)
         );
  AOI22_X1 U73 ( .A1(n194), .A2(n140), .B1(LU_OpA[21]), .B2(n200), .ZN(n139)
         );
  AOI22_X1 U74 ( .A1(n194), .A2(n136), .B1(LU_OpA[22]), .B2(n200), .ZN(n135)
         );
  AOI22_X1 U75 ( .A1(n194), .A2(n132), .B1(LU_OpA[23]), .B2(n200), .ZN(n131)
         );
  AOI22_X1 U76 ( .A1(n193), .A2(n156), .B1(LU_OpA[18]), .B2(n199), .ZN(n155)
         );
  AOI22_X1 U77 ( .A1(n193), .A2(n152), .B1(LU_OpA[19]), .B2(n199), .ZN(n151)
         );
  AOI22_X1 U78 ( .A1(n193), .A2(n160), .B1(LU_OpA[17]), .B2(n199), .ZN(n159)
         );
  AOI22_X1 U79 ( .A1(n193), .A2(n148), .B1(LU_OpA[1]), .B2(n199), .ZN(n147) );
  AOI22_X1 U80 ( .A1(n193), .A2(n172), .B1(LU_OpA[14]), .B2(n199), .ZN(n171)
         );
  AOI22_X1 U81 ( .A1(n193), .A2(n176), .B1(LU_OpA[13]), .B2(n199), .ZN(n175)
         );
  AOI22_X1 U82 ( .A1(n193), .A2(n168), .B1(LU_OpA[15]), .B2(n199), .ZN(n167)
         );
  AOI22_X1 U83 ( .A1(n193), .A2(n164), .B1(LU_OpA[16]), .B2(n199), .ZN(n163)
         );
  AOI22_X1 U84 ( .A1(n194), .A2(n112), .B1(LU_OpA[28]), .B2(n200), .ZN(n111)
         );
  AOI22_X1 U85 ( .A1(n194), .A2(n108), .B1(LU_OpA[29]), .B2(n200), .ZN(n107)
         );
  AOI22_X1 U86 ( .A1(n194), .A2(n104), .B1(LU_OpA[2]), .B2(n200), .ZN(n103) );
  AOI22_X1 U87 ( .A1(n194), .A2(n128), .B1(LU_OpA[24]), .B2(n200), .ZN(n127)
         );
  AOI22_X1 U88 ( .A1(n194), .A2(n120), .B1(LU_OpA[26]), .B2(n200), .ZN(n119)
         );
  AOI22_X1 U89 ( .A1(n194), .A2(n124), .B1(LU_OpA[25]), .B2(n200), .ZN(n123)
         );
  AOI22_X1 U90 ( .A1(n194), .A2(n116), .B1(LU_OpA[27]), .B2(n200), .ZN(n115)
         );
  AOI22_X1 U91 ( .A1(n198), .A2(n92), .B1(LU_OpA[3]), .B2(n204), .ZN(n89) );
  AOI22_X1 U92 ( .A1(n198), .A2(n88), .B1(LU_OpA[4]), .B2(n204), .ZN(n85) );
  AOI22_X1 U93 ( .A1(n198), .A2(n84), .B1(LU_OpA[5]), .B2(n204), .ZN(n81) );
  AOI22_X1 U94 ( .A1(n198), .A2(n72), .B1(LU_OpA[8]), .B2(n204), .ZN(n69) );
  AOI22_X1 U95 ( .A1(n198), .A2(n76), .B1(LU_OpA[7]), .B2(n204), .ZN(n73) );
  AOI22_X1 U96 ( .A1(n198), .A2(n80), .B1(LU_OpA[6]), .B2(n204), .ZN(n77) );
  AOI22_X1 U97 ( .A1(n198), .A2(n68), .B1(n204), .B2(LU_OpA[9]), .ZN(n65) );
  AOI22_X1 U98 ( .A1(n196), .A2(n192), .B1(LU_OpA[0]), .B2(n202), .ZN(n189) );
  AOI22_X1 U99 ( .A1(n196), .A2(n180), .B1(LU_OpA[12]), .B2(n202), .ZN(n177)
         );
  AOI22_X1 U100 ( .A1(n196), .A2(n188), .B1(LU_OpA[10]), .B2(n202), .ZN(n185)
         );
  AOI22_X1 U101 ( .A1(n196), .A2(n184), .B1(LU_OpA[11]), .B2(n202), .ZN(n181)
         );
  AOI22_X1 U102 ( .A1(n197), .A2(n144), .B1(LU_OpA[20]), .B2(n203), .ZN(n141)
         );
  AOI22_X1 U103 ( .A1(n197), .A2(n140), .B1(LU_OpA[21]), .B2(n203), .ZN(n137)
         );
  AOI22_X1 U104 ( .A1(n197), .A2(n136), .B1(LU_OpA[22]), .B2(n203), .ZN(n133)
         );
  AOI22_X1 U105 ( .A1(n197), .A2(n132), .B1(LU_OpA[23]), .B2(n203), .ZN(n129)
         );
  AOI22_X1 U106 ( .A1(n196), .A2(n156), .B1(LU_OpA[18]), .B2(n202), .ZN(n153)
         );
  AOI22_X1 U107 ( .A1(n196), .A2(n152), .B1(LU_OpA[19]), .B2(n202), .ZN(n149)
         );
  AOI22_X1 U108 ( .A1(n196), .A2(n160), .B1(LU_OpA[17]), .B2(n202), .ZN(n157)
         );
  AOI22_X1 U109 ( .A1(n196), .A2(n148), .B1(LU_OpA[1]), .B2(n202), .ZN(n145)
         );
  AOI22_X1 U110 ( .A1(n196), .A2(n172), .B1(LU_OpA[14]), .B2(n202), .ZN(n169)
         );
  AOI22_X1 U111 ( .A1(n196), .A2(n176), .B1(LU_OpA[13]), .B2(n202), .ZN(n173)
         );
  AOI22_X1 U112 ( .A1(n196), .A2(n168), .B1(LU_OpA[15]), .B2(n202), .ZN(n165)
         );
  AOI22_X1 U113 ( .A1(n196), .A2(n164), .B1(LU_OpA[16]), .B2(n202), .ZN(n161)
         );
  AOI22_X1 U114 ( .A1(n197), .A2(n112), .B1(LU_OpA[28]), .B2(n203), .ZN(n109)
         );
  AOI22_X1 U115 ( .A1(n197), .A2(n108), .B1(LU_OpA[29]), .B2(n203), .ZN(n105)
         );
  AOI22_X1 U116 ( .A1(n197), .A2(n104), .B1(LU_OpA[2]), .B2(n203), .ZN(n101)
         );
  AOI22_X1 U117 ( .A1(n197), .A2(n128), .B1(LU_OpA[24]), .B2(n203), .ZN(n125)
         );
  AOI22_X1 U118 ( .A1(n197), .A2(n120), .B1(LU_OpA[26]), .B2(n203), .ZN(n117)
         );
  AOI22_X1 U119 ( .A1(n197), .A2(n124), .B1(LU_OpA[25]), .B2(n203), .ZN(n121)
         );
  AOI22_X1 U120 ( .A1(n197), .A2(n116), .B1(LU_OpA[27]), .B2(n203), .ZN(n113)
         );
  OAI22_X1 U121 ( .A1(n101), .A2(n102), .B1(LU_OpB[2]), .B2(n103), .ZN(LU_Y[2]) );
  INV_X1 U122 ( .A(LU_OpB[2]), .ZN(n102) );
  BUF_X1 U123 ( .A(LU_Opcode[1]), .Z(n196) );
  BUF_X1 U124 ( .A(LU_Opcode[1]), .Z(n197) );
  BUF_X1 U125 ( .A(LU_Opcode[1]), .Z(n198) );
  OAI22_X1 U126 ( .A1(n137), .A2(n138), .B1(LU_OpB[21]), .B2(n139), .ZN(
        LU_Y[21]) );
  INV_X1 U127 ( .A(LU_OpB[21]), .ZN(n138) );
  OAI22_X1 U128 ( .A1(n157), .A2(n158), .B1(LU_OpB[17]), .B2(n159), .ZN(
        LU_Y[17]) );
  INV_X1 U129 ( .A(LU_OpB[17]), .ZN(n158) );
  OAI22_X1 U130 ( .A1(n173), .A2(n174), .B1(LU_OpB[13]), .B2(n175), .ZN(
        LU_Y[13]) );
  INV_X1 U131 ( .A(LU_OpB[13]), .ZN(n174) );
  OAI22_X1 U132 ( .A1(n105), .A2(n106), .B1(LU_OpB[29]), .B2(n107), .ZN(
        LU_Y[29]) );
  INV_X1 U133 ( .A(LU_OpB[29]), .ZN(n106) );
  OAI22_X1 U134 ( .A1(n121), .A2(n122), .B1(LU_OpB[25]), .B2(n123), .ZN(
        LU_Y[25]) );
  INV_X1 U135 ( .A(LU_OpB[25]), .ZN(n122) );
  OAI22_X1 U136 ( .A1(n65), .A2(n66), .B1(LU_OpB[9]), .B2(n67), .ZN(LU_Y[9])
         );
  INV_X1 U137 ( .A(LU_OpB[9]), .ZN(n66) );
  OAI22_X1 U138 ( .A1(n81), .A2(n82), .B1(LU_OpB[5]), .B2(n83), .ZN(LU_Y[5])
         );
  INV_X1 U139 ( .A(LU_OpB[5]), .ZN(n82) );
  OAI22_X1 U140 ( .A1(n145), .A2(n146), .B1(LU_OpB[1]), .B2(n147), .ZN(LU_Y[1]) );
  INV_X1 U141 ( .A(LU_OpB[1]), .ZN(n146) );
  BUF_X1 U142 ( .A(LU_Opcode[0]), .Z(n193) );
  BUF_X1 U143 ( .A(LU_Opcode[0]), .Z(n194) );
  BUF_X1 U144 ( .A(LU_Opcode[2]), .Z(n199) );
  BUF_X1 U145 ( .A(LU_Opcode[3]), .Z(n202) );
  BUF_X1 U146 ( .A(LU_Opcode[2]), .Z(n200) );
  BUF_X1 U147 ( .A(LU_Opcode[3]), .Z(n203) );
  BUF_X1 U148 ( .A(LU_Opcode[2]), .Z(n201) );
  BUF_X1 U149 ( .A(LU_Opcode[3]), .Z(n204) );
  BUF_X1 U150 ( .A(LU_Opcode[0]), .Z(n195) );
  OAI22_X1 U151 ( .A1(n177), .A2(n178), .B1(LU_OpB[12]), .B2(n179), .ZN(
        LU_Y[12]) );
  INV_X1 U152 ( .A(LU_OpB[12]), .ZN(n178) );
  OAI22_X1 U153 ( .A1(n141), .A2(n142), .B1(LU_OpB[20]), .B2(n143), .ZN(
        LU_Y[20]) );
  INV_X1 U154 ( .A(LU_OpB[20]), .ZN(n142) );
  OAI22_X1 U155 ( .A1(n161), .A2(n162), .B1(LU_OpB[16]), .B2(n163), .ZN(
        LU_Y[16]) );
  INV_X1 U156 ( .A(LU_OpB[16]), .ZN(n162) );
  OAI22_X1 U157 ( .A1(n109), .A2(n110), .B1(LU_OpB[28]), .B2(n111), .ZN(
        LU_Y[28]) );
  INV_X1 U158 ( .A(LU_OpB[28]), .ZN(n110) );
  OAI22_X1 U159 ( .A1(n125), .A2(n126), .B1(LU_OpB[24]), .B2(n127), .ZN(
        LU_Y[24]) );
  INV_X1 U160 ( .A(LU_OpB[24]), .ZN(n126) );
  OAI22_X1 U161 ( .A1(n69), .A2(n70), .B1(LU_OpB[8]), .B2(n71), .ZN(LU_Y[8])
         );
  INV_X1 U162 ( .A(LU_OpB[8]), .ZN(n70) );
  OAI22_X1 U163 ( .A1(n85), .A2(n86), .B1(LU_OpB[4]), .B2(n87), .ZN(LU_Y[4])
         );
  INV_X1 U164 ( .A(LU_OpB[4]), .ZN(n86) );
  OAI22_X1 U165 ( .A1(n189), .A2(n190), .B1(LU_OpB[0]), .B2(n191), .ZN(LU_Y[0]) );
  INV_X1 U166 ( .A(LU_OpB[0]), .ZN(n190) );
  AOI22_X1 U167 ( .A1(n197), .A2(n100), .B1(LU_OpA[30]), .B2(n203), .ZN(n97)
         );
  AOI22_X1 U168 ( .A1(n194), .A2(n100), .B1(LU_OpA[30]), .B2(n200), .ZN(n99)
         );
  INV_X1 U169 ( .A(LU_OpA[30]), .ZN(n100) );
  AOI22_X1 U170 ( .A1(n198), .A2(n96), .B1(LU_OpA[31]), .B2(n204), .ZN(n93) );
  AOI22_X1 U171 ( .A1(n195), .A2(n96), .B1(LU_OpA[31]), .B2(n201), .ZN(n95) );
  INV_X1 U172 ( .A(LU_OpA[31]), .ZN(n96) );
endmodule


module P4Adder_N32 ( A, B, c_in, c_out, Sum );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Sum;
  input c_in;
  output c_out;

  wire   [7:1] carry_tmp;

  CarryGenerator_N32_K8 CG ( .A(A), .B(B), .c_in(c_in), .CarryVector({c_out, 
        carry_tmp}) );
  CarrySelect_N32_K4 CS ( .A(A), .B(B), .Cin({carry_tmp, c_in}), .S(Sum) );
endmodule


module Barrel_Shifter_NBIT_AMOUNT5 ( BS_data_in, BS_opcode, BS_amount, 
        BS_data_out );
  input [31:0] BS_data_in;
  input [1:0] BS_opcode;
  input [4:0] BS_amount;
  output [31:0] BS_data_out;
  wire   \s_mX2[0][0][39] , \s_mX2[0][0][38] , \s_mX2[0][0][37] ,
         \s_mX2[0][0][36] , \s_mX2[0][0][35] , \s_mX2[0][0][34] ,
         \s_mX2[0][0][33] , \s_mX2[0][0][32] , \s_mX2[0][0][31] ,
         \s_mX2[0][0][30] , \s_mX2[0][0][29] , \s_mX2[0][0][28] ,
         \s_mX2[0][0][27] , \s_mX2[0][0][26] , \s_mX2[0][0][25] ,
         \s_mX2[0][0][24] , \s_mX2[0][0][23] , \s_mX2[0][0][22] ,
         \s_mX2[0][0][21] , \s_mX2[0][0][20] , \s_mX2[0][0][19] ,
         \s_mX2[0][0][18] , \s_mX2[0][0][17] , \s_mX2[0][0][16] ,
         \s_mX2[0][0][15] , \s_mX2[0][0][14] , \s_mX2[0][0][13] ,
         \s_mX2[0][0][12] , \s_mX2[0][0][11] , \s_mX2[0][0][10] ,
         \s_mX2[0][0][9] , \s_mX2[0][0][8] , \s_mX2[0][0][7] ,
         \s_mX2[0][0][6] , \s_mX2[0][0][5] , \s_mX2[0][0][4] ,
         \s_mX2[0][0][3] , \s_mX2[0][0][2] , \s_mX2[0][0][1] ,
         \s_mX2[0][0][0] , \s_mX2[0][1][39] , \s_mX2[0][1][38] ,
         \s_mX2[0][1][37] , \s_mX2[0][1][36] , \s_mX2[0][1][35] ,
         \s_mX2[0][1][34] , \s_mX2[0][1][33] , \s_mX2[0][1][32] ,
         \s_mX2[0][1][31] , \s_mX2[0][1][30] , \s_mX2[0][1][29] ,
         \s_mX2[0][1][28] , \s_mX2[0][1][27] , \s_mX2[0][1][26] ,
         \s_mX2[0][1][25] , \s_mX2[0][1][24] , \s_mX2[0][1][23] ,
         \s_mX2[0][1][22] , \s_mX2[0][1][21] , \s_mX2[0][1][20] ,
         \s_mX2[0][1][19] , \s_mX2[0][1][18] , \s_mX2[0][1][17] ,
         \s_mX2[0][1][16] , \s_mX2[0][1][15] , \s_mX2[0][1][14] ,
         \s_mX2[0][1][13] , \s_mX2[0][1][12] , \s_mX2[0][1][11] ,
         \s_mX2[0][1][10] , \s_mX2[0][1][9] , \s_mX2[0][1][8] ,
         \s_mX2[0][1][7] , \s_mX2[0][1][6] , \s_mX2[0][1][5] ,
         \s_mX2[0][1][4] , \s_mX2[0][1][3] , \s_mX2[0][1][2] ,
         \s_mX2[0][1][1] , \s_mX2[0][1][0] , \s_mX2[0][2][39] ,
         \s_mX2[0][2][38] , \s_mX2[0][2][37] , \s_mX2[0][2][36] ,
         \s_mX2[0][2][35] , \s_mX2[0][2][34] , \s_mX2[0][2][33] ,
         \s_mX2[0][2][32] , \s_mX2[0][2][31] , \s_mX2[0][2][30] ,
         \s_mX2[0][2][29] , \s_mX2[0][2][28] , \s_mX2[0][2][27] ,
         \s_mX2[0][2][26] , \s_mX2[0][2][25] , \s_mX2[0][2][24] ,
         \s_mX2[0][2][23] , \s_mX2[0][2][22] , \s_mX2[0][2][21] ,
         \s_mX2[0][2][20] , \s_mX2[0][2][19] , \s_mX2[0][2][18] ,
         \s_mX2[0][2][17] , \s_mX2[0][2][16] , \s_mX2[0][2][15] ,
         \s_mX2[0][2][14] , \s_mX2[0][2][13] , \s_mX2[0][2][12] ,
         \s_mX2[0][2][11] , \s_mX2[0][2][10] , \s_mX2[0][2][9] ,
         \s_mX2[0][2][8] , \s_mX2[0][2][7] , \s_mX2[0][2][6] ,
         \s_mX2[0][2][5] , \s_mX2[0][2][4] , \s_mX2[0][2][3] ,
         \s_mX2[0][2][2] , \s_mX2[0][2][1] , \s_mX2[0][2][0] ,
         \s_mX2[0][3][39] , \s_mX2[0][3][38] , \s_mX2[0][3][37] ,
         \s_mX2[0][3][36] , \s_mX2[0][3][35] , \s_mX2[0][3][34] ,
         \s_mX2[0][3][33] , \s_mX2[0][3][32] , \s_mX2[0][3][31] ,
         \s_mX2[0][3][30] , \s_mX2[0][3][29] , \s_mX2[0][3][28] ,
         \s_mX2[0][3][27] , \s_mX2[0][3][26] , \s_mX2[0][3][25] ,
         \s_mX2[0][3][24] , \s_mX2[0][3][23] , \s_mX2[0][3][22] ,
         \s_mX2[0][3][21] , \s_mX2[0][3][20] , \s_mX2[0][3][19] ,
         \s_mX2[0][3][18] , \s_mX2[0][3][17] , \s_mX2[0][3][16] ,
         \s_mX2[0][3][15] , \s_mX2[0][3][14] , \s_mX2[0][3][13] ,
         \s_mX2[0][3][12] , \s_mX2[0][3][11] , \s_mX2[0][3][10] ,
         \s_mX2[0][3][9] , \s_mX2[0][3][8] , \s_mX2[0][3][7] ,
         \s_mX2[0][3][6] , \s_mX2[0][3][5] , \s_mX2[0][3][4] ,
         \s_mX2[0][3][3] , \s_mX2[0][3][2] , \s_mX2[0][3][1] ,
         \s_mX2[0][3][0] , \s_mX2[1][0][39] , \s_mX2[1][0][38] ,
         \s_mX2[1][0][37] , \s_mX2[1][0][36] , \s_mX2[1][0][35] ,
         \s_mX2[1][0][34] , \s_mX2[1][0][33] , \s_mX2[1][0][32] ,
         \s_mX2[1][0][31] , \s_mX2[1][0][30] , \s_mX2[1][0][29] ,
         \s_mX2[1][0][28] , \s_mX2[1][0][27] , \s_mX2[1][0][26] ,
         \s_mX2[1][0][25] , \s_mX2[1][0][24] , \s_mX2[1][0][23] ,
         \s_mX2[1][0][22] , \s_mX2[1][0][21] , \s_mX2[1][0][20] ,
         \s_mX2[1][0][19] , \s_mX2[1][0][18] , \s_mX2[1][0][17] ,
         \s_mX2[1][0][16] , \s_mX2[1][0][15] , \s_mX2[1][0][14] ,
         \s_mX2[1][0][13] , \s_mX2[1][0][12] , \s_mX2[1][0][11] ,
         \s_mX2[1][0][10] , \s_mX2[1][0][9] , \s_mX2[1][0][8] ,
         \s_mX2[1][0][7] , \s_mX2[1][0][6] , \s_mX2[1][0][5] ,
         \s_mX2[1][0][4] , \s_mX2[1][0][3] , \s_mX2[1][0][2] ,
         \s_mX2[1][0][1] , \s_mX2[1][0][0] , \s_mX2[1][2][39] ,
         \s_mX2[1][2][38] , \s_mX2[1][2][37] , \s_mX2[1][2][36] ,
         \s_mX2[1][2][35] , \s_mX2[1][2][34] , \s_mX2[1][2][33] ,
         \s_mX2[1][2][32] , \s_mX2[1][2][31] , \s_mX2[1][2][30] ,
         \s_mX2[1][2][29] , \s_mX2[1][2][28] , \s_mX2[1][2][27] ,
         \s_mX2[1][2][26] , \s_mX2[1][2][25] , \s_mX2[1][2][24] ,
         \s_mX2[1][2][23] , \s_mX2[1][2][22] , \s_mX2[1][2][21] ,
         \s_mX2[1][2][20] , \s_mX2[1][2][19] , \s_mX2[1][2][18] ,
         \s_mX2[1][2][17] , \s_mX2[1][2][16] , \s_mX2[1][2][15] ,
         \s_mX2[1][2][14] , \s_mX2[1][2][13] , \s_mX2[1][2][12] ,
         \s_mX2[1][2][11] , \s_mX2[1][2][10] , \s_mX2[1][2][9] ,
         \s_mX2[1][2][8] , \s_mX2[1][2][7] , \s_mX2[1][2][6] ,
         \s_mX2[1][2][5] , \s_mX2[1][2][4] , \s_mX2[1][2][3] ,
         \s_mX2[1][2][2] , \s_mX2[1][2][1] , \s_mX2[1][2][0] ,
         \s_mX2[2][0][39] , \s_mX2[2][0][38] , \s_mX2[2][0][37] ,
         \s_mX2[2][0][36] , \s_mX2[2][0][35] , \s_mX2[2][0][34] ,
         \s_mX2[2][0][33] , \s_mX2[2][0][32] , \s_mX2[2][0][31] ,
         \s_mX2[2][0][30] , \s_mX2[2][0][29] , \s_mX2[2][0][28] ,
         \s_mX2[2][0][27] , \s_mX2[2][0][26] , \s_mX2[2][0][25] ,
         \s_mX2[2][0][24] , \s_mX2[2][0][23] , \s_mX2[2][0][22] ,
         \s_mX2[2][0][21] , \s_mX2[2][0][20] , \s_mX2[2][0][19] ,
         \s_mX2[2][0][18] , \s_mX2[2][0][17] , \s_mX2[2][0][16] ,
         \s_mX2[2][0][15] , \s_mX2[2][0][14] , \s_mX2[2][0][13] ,
         \s_mX2[2][0][12] , \s_mX2[2][0][11] , \s_mX2[2][0][10] ,
         \s_mX2[2][0][9] , \s_mX2[2][0][8] , \s_mX2[2][0][7] ,
         \s_mX2[2][0][6] , \s_mX2[2][0][5] , \s_mX2[2][0][4] ,
         \s_mX2[2][0][3] , \s_mX2[2][0][2] , \s_mX2[2][0][1] ,
         \s_mX2[2][0][0] , \s_out_mask[1][0][31] , \s_out_mask[1][0][30] ,
         \s_out_mask[1][0][29] , \s_out_mask[1][0][28] ,
         \s_out_mask[1][0][27] , \s_out_mask[1][0][26] ,
         \s_out_mask[1][0][25] , \s_out_mask[1][0][24] ,
         \s_out_mask[1][0][23] , \s_out_mask[1][0][22] ,
         \s_out_mask[1][0][21] , \s_out_mask[1][0][20] ,
         \s_out_mask[1][0][19] , \s_out_mask[1][0][18] ,
         \s_out_mask[1][0][17] , \s_out_mask[1][0][16] ,
         \s_out_mask[1][0][15] , \s_out_mask[1][0][14] ,
         \s_out_mask[1][0][13] , \s_out_mask[1][0][12] ,
         \s_out_mask[1][0][11] , \s_out_mask[1][0][10] , \s_out_mask[1][0][9] ,
         \s_out_mask[1][0][8] , \s_out_mask[1][0][7] , \s_out_mask[1][0][6] ,
         \s_out_mask[1][0][5] , \s_out_mask[1][0][4] , \s_out_mask[1][0][3] ,
         \s_out_mask[1][0][2] , \s_out_mask[1][0][1] , \s_out_mask[1][0][0] ,
         \s_out_mask[1][2][31] , \s_out_mask[1][2][30] ,
         \s_out_mask[1][2][29] , \s_out_mask[1][2][28] ,
         \s_out_mask[1][2][27] , \s_out_mask[1][2][26] ,
         \s_out_mask[1][2][25] , \s_out_mask[1][2][24] ,
         \s_out_mask[1][2][23] , \s_out_mask[1][2][22] ,
         \s_out_mask[1][2][21] , \s_out_mask[1][2][20] ,
         \s_out_mask[1][2][19] , \s_out_mask[1][2][18] ,
         \s_out_mask[1][2][17] , \s_out_mask[1][2][16] ,
         \s_out_mask[1][2][15] , \s_out_mask[1][2][14] ,
         \s_out_mask[1][2][13] , \s_out_mask[1][2][12] ,
         \s_out_mask[1][2][11] , \s_out_mask[1][2][10] , \s_out_mask[1][2][9] ,
         \s_out_mask[1][2][8] , \s_out_mask[1][2][7] , \s_out_mask[1][2][6] ,
         \s_out_mask[1][2][5] , \s_out_mask[1][2][4] , \s_out_mask[1][2][3] ,
         \s_out_mask[1][2][2] , \s_out_mask[1][2][1] , \s_out_mask[1][2][0] ,
         \s_out_mask[1][4][31] , \s_out_mask[1][4][30] ,
         \s_out_mask[1][4][29] , \s_out_mask[1][4][28] ,
         \s_out_mask[1][4][27] , \s_out_mask[1][4][26] ,
         \s_out_mask[1][4][25] , \s_out_mask[1][4][24] ,
         \s_out_mask[1][4][23] , \s_out_mask[1][4][22] ,
         \s_out_mask[1][4][21] , \s_out_mask[1][4][20] ,
         \s_out_mask[1][4][19] , \s_out_mask[1][4][18] ,
         \s_out_mask[1][4][17] , \s_out_mask[1][4][16] ,
         \s_out_mask[1][4][15] , \s_out_mask[1][4][14] ,
         \s_out_mask[1][4][13] , \s_out_mask[1][4][12] ,
         \s_out_mask[1][4][11] , \s_out_mask[1][4][10] , \s_out_mask[1][4][9] ,
         \s_out_mask[1][4][8] , \s_out_mask[1][4][7] , \s_out_mask[1][4][6] ,
         \s_out_mask[1][4][5] , \s_out_mask[1][4][4] , \s_out_mask[1][4][3] ,
         \s_out_mask[1][4][2] , \s_out_mask[1][4][1] , \s_out_mask[1][4][0] ,
         \s_out_mask[1][6][31] , \s_out_mask[1][6][30] ,
         \s_out_mask[1][6][29] , \s_out_mask[1][6][28] ,
         \s_out_mask[1][6][27] , \s_out_mask[1][6][26] ,
         \s_out_mask[1][6][25] , \s_out_mask[1][6][24] ,
         \s_out_mask[1][6][23] , \s_out_mask[1][6][22] ,
         \s_out_mask[1][6][21] , \s_out_mask[1][6][20] ,
         \s_out_mask[1][6][19] , \s_out_mask[1][6][18] ,
         \s_out_mask[1][6][17] , \s_out_mask[1][6][16] ,
         \s_out_mask[1][6][15] , \s_out_mask[1][6][14] ,
         \s_out_mask[1][6][13] , \s_out_mask[1][6][12] ,
         \s_out_mask[1][6][11] , \s_out_mask[1][6][10] , \s_out_mask[1][6][9] ,
         \s_out_mask[1][6][8] , \s_out_mask[1][6][7] , \s_out_mask[1][6][6] ,
         \s_out_mask[1][6][5] , \s_out_mask[1][6][4] , \s_out_mask[1][6][3] ,
         \s_out_mask[1][6][2] , \s_out_mask[1][6][1] , \s_out_mask[1][6][0] ,
         \s_out_mask[2][0][31] , \s_out_mask[2][0][30] ,
         \s_out_mask[2][0][29] , \s_out_mask[2][0][28] ,
         \s_out_mask[2][0][27] , \s_out_mask[2][0][26] ,
         \s_out_mask[2][0][25] , \s_out_mask[2][0][24] ,
         \s_out_mask[2][0][23] , \s_out_mask[2][0][22] ,
         \s_out_mask[2][0][21] , \s_out_mask[2][0][20] ,
         \s_out_mask[2][0][19] , \s_out_mask[2][0][18] ,
         \s_out_mask[2][0][17] , \s_out_mask[2][0][16] ,
         \s_out_mask[2][0][15] , \s_out_mask[2][0][14] ,
         \s_out_mask[2][0][13] , \s_out_mask[2][0][12] ,
         \s_out_mask[2][0][11] , \s_out_mask[2][0][10] , \s_out_mask[2][0][9] ,
         \s_out_mask[2][0][8] , \s_out_mask[2][0][7] , \s_out_mask[2][0][6] ,
         \s_out_mask[2][0][5] , \s_out_mask[2][0][4] , \s_out_mask[2][0][3] ,
         \s_out_mask[2][0][2] , \s_out_mask[2][0][1] , \s_out_mask[2][0][0] ,
         \s_out_mask[2][4][31] , \s_out_mask[2][4][30] ,
         \s_out_mask[2][4][29] , \s_out_mask[2][4][28] ,
         \s_out_mask[2][4][27] , \s_out_mask[2][4][26] ,
         \s_out_mask[2][4][25] , \s_out_mask[2][4][24] ,
         \s_out_mask[2][4][23] , \s_out_mask[2][4][22] ,
         \s_out_mask[2][4][21] , \s_out_mask[2][4][20] ,
         \s_out_mask[2][4][19] , \s_out_mask[2][4][18] ,
         \s_out_mask[2][4][17] , \s_out_mask[2][4][16] ,
         \s_out_mask[2][4][15] , \s_out_mask[2][4][14] ,
         \s_out_mask[2][4][13] , \s_out_mask[2][4][12] ,
         \s_out_mask[2][4][11] , \s_out_mask[2][4][10] , \s_out_mask[2][4][9] ,
         \s_out_mask[2][4][8] , \s_out_mask[2][4][7] , \s_out_mask[2][4][6] ,
         \s_out_mask[2][4][5] , \s_out_mask[2][4][4] , \s_out_mask[2][4][3] ,
         \s_out_mask[2][4][2] , \s_out_mask[2][4][1] , \s_out_mask[2][4][0] ,
         n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18,
         n19, n20, n21, n22, n23, n24, n25, n26;
  wire   [7:0] s_msb;
  wire   [39:1] s_selected_mask;
  wire   [2:0] s_amount;
  wire   [2:0] s_not_amount;
  wire   [2:0] s_sel_out;
  wire   SYNOPSYS_UNCONNECTED__0;
  assign n4 = BS_opcode[0];

  Mux_NBit_2x1_NBIT_IN8_0 MSB_MUX ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0}), .port1({BS_data_in[31], BS_data_in[31], BS_data_in[31], 
        BS_data_in[31], BS_data_in[31], BS_data_in[31], BS_data_in[31], 
        BS_data_in[31]}), .sel(BS_opcode[1]), .portY(s_msb) );
  Mux_NBit_2x1_NBIT_IN8_20 MUX2_0_0 ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .port1(BS_data_in[7:0]), .sel(n23), .portY({
        \s_mX2[0][0][7] , \s_mX2[0][0][6] , \s_mX2[0][0][5] , \s_mX2[0][0][4] , 
        \s_mX2[0][0][3] , \s_mX2[0][0][2] , \s_mX2[0][0][1] , \s_mX2[0][0][0] }) );
  Mux_NBit_2x1_NBIT_IN8_19 MUX1_0_1 ( .port0(BS_data_in[7:0]), .port1(
        BS_data_in[15:8]), .sel(n26), .portY({\s_mX2[0][0][15] , 
        \s_mX2[0][0][14] , \s_mX2[0][0][13] , \s_mX2[0][0][12] , 
        \s_mX2[0][0][11] , \s_mX2[0][0][10] , \s_mX2[0][0][9] , 
        \s_mX2[0][0][8] }) );
  Mux_NBit_2x1_NBIT_IN8_18 MUX1_0_2 ( .port0(BS_data_in[15:8]), .port1(
        BS_data_in[23:16]), .sel(n26), .portY({\s_mX2[0][0][23] , 
        \s_mX2[0][0][22] , \s_mX2[0][0][21] , \s_mX2[0][0][20] , 
        \s_mX2[0][0][19] , \s_mX2[0][0][18] , \s_mX2[0][0][17] , 
        \s_mX2[0][0][16] }) );
  Mux_NBit_2x1_NBIT_IN8_17 MUX1_0_3 ( .port0(BS_data_in[23:16]), .port1(
        BS_data_in[31:24]), .sel(n25), .portY({\s_mX2[0][0][31] , 
        \s_mX2[0][0][30] , \s_mX2[0][0][29] , \s_mX2[0][0][28] , 
        \s_mX2[0][0][27] , \s_mX2[0][0][26] , \s_mX2[0][0][25] , 
        \s_mX2[0][0][24] }) );
  Mux_NBit_2x1_NBIT_IN8_16 MUX3_0_4 ( .port0({n10, BS_data_in[30:24]}), 
        .port1(s_msb), .sel(n25), .portY({\s_mX2[0][0][39] , \s_mX2[0][0][38] , 
        \s_mX2[0][0][37] , \s_mX2[0][0][36] , \s_mX2[0][0][35] , 
        \s_mX2[0][0][34] , \s_mX2[0][0][33] , \s_mX2[0][0][32] }) );
  Mux_NBit_2x1_NBIT_IN8_15 MUX2_1_0 ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .port1(BS_data_in[15:8]), .sel(n25), .portY({
        \s_mX2[0][1][7] , \s_mX2[0][1][6] , \s_mX2[0][1][5] , \s_mX2[0][1][4] , 
        \s_mX2[0][1][3] , \s_mX2[0][1][2] , \s_mX2[0][1][1] , \s_mX2[0][1][0] }) );
  Mux_NBit_2x1_NBIT_IN8_14 MUX2_1_1 ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .port1(BS_data_in[23:16]), .sel(n24), .portY({
        \s_mX2[0][1][15] , \s_mX2[0][1][14] , \s_mX2[0][1][13] , 
        \s_mX2[0][1][12] , \s_mX2[0][1][11] , \s_mX2[0][1][10] , 
        \s_mX2[0][1][9] , \s_mX2[0][1][8] }) );
  Mux_NBit_2x1_NBIT_IN8_13 MUX1_1_2 ( .port0(BS_data_in[7:0]), .port1({n10, 
        BS_data_in[30:24]}), .sel(n24), .portY({\s_mX2[0][1][23] , 
        \s_mX2[0][1][22] , \s_mX2[0][1][21] , \s_mX2[0][1][20] , 
        \s_mX2[0][1][19] , \s_mX2[0][1][18] , \s_mX2[0][1][17] , 
        \s_mX2[0][1][16] }) );
  Mux_NBit_2x1_NBIT_IN8_12 MUX3_1_3 ( .port0(BS_data_in[15:8]), .port1(s_msb), 
        .sel(n24), .portY({\s_mX2[0][1][31] , \s_mX2[0][1][30] , 
        \s_mX2[0][1][29] , \s_mX2[0][1][28] , \s_mX2[0][1][27] , 
        \s_mX2[0][1][26] , \s_mX2[0][1][25] , \s_mX2[0][1][24] }) );
  Mux_NBit_2x1_NBIT_IN8_11 MUX3_1_4 ( .port0(BS_data_in[23:16]), .port1(s_msb), 
        .sel(n23), .portY({\s_mX2[0][1][39] , \s_mX2[0][1][38] , 
        \s_mX2[0][1][37] , \s_mX2[0][1][36] , \s_mX2[0][1][35] , 
        \s_mX2[0][1][34] , \s_mX2[0][1][33] , \s_mX2[0][1][32] }) );
  Mux_NBit_2x1_NBIT_IN8_10 MUX2_2_0 ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .port1(BS_data_in[23:16]), .sel(n23), .portY({
        \s_mX2[0][2][7] , \s_mX2[0][2][6] , \s_mX2[0][2][5] , \s_mX2[0][2][4] , 
        \s_mX2[0][2][3] , \s_mX2[0][2][2] , \s_mX2[0][2][1] , \s_mX2[0][2][0] }) );
  Mux_NBit_2x1_NBIT_IN8_9 MUX2_2_1 ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .port1({n10, BS_data_in[30:24]}), .sel(n22), 
        .portY({\s_mX2[0][2][15] , \s_mX2[0][2][14] , \s_mX2[0][2][13] , 
        \s_mX2[0][2][12] , \s_mX2[0][2][11] , \s_mX2[0][2][10] , 
        \s_mX2[0][2][9] , \s_mX2[0][2][8] }) );
  Mux_NBit_2x1_NBIT_IN8_8 MUX4_2_2 ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .port1({s_msb[7:3], n7, s_msb[1], n8}), .sel(n22), 
        .portY({\s_mX2[0][2][23] , \s_mX2[0][2][22] , \s_mX2[0][2][21] , 
        \s_mX2[0][2][20] , \s_mX2[0][2][19] , \s_mX2[0][2][18] , 
        \s_mX2[0][2][17] , \s_mX2[0][2][16] }) );
  Mux_NBit_2x1_NBIT_IN8_7 MUX3_2_3 ( .port0(BS_data_in[7:0]), .port1(s_msb), 
        .sel(n22), .portY({\s_mX2[0][2][31] , \s_mX2[0][2][30] , 
        \s_mX2[0][2][29] , \s_mX2[0][2][28] , \s_mX2[0][2][27] , 
        \s_mX2[0][2][26] , \s_mX2[0][2][25] , \s_mX2[0][2][24] }) );
  Mux_NBit_2x1_NBIT_IN8_6 MUX3_2_4 ( .port0(BS_data_in[15:8]), .port1(s_msb), 
        .sel(n21), .portY({\s_mX2[0][2][39] , \s_mX2[0][2][38] , 
        \s_mX2[0][2][37] , \s_mX2[0][2][36] , \s_mX2[0][2][35] , 
        \s_mX2[0][2][34] , \s_mX2[0][2][33] , \s_mX2[0][2][32] }) );
  Mux_NBit_2x1_NBIT_IN8_5 MUX2_3_0 ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .port1({n10, BS_data_in[30:24]}), .sel(n21), 
        .portY({\s_mX2[0][3][7] , \s_mX2[0][3][6] , \s_mX2[0][3][5] , 
        \s_mX2[0][3][4] , \s_mX2[0][3][3] , \s_mX2[0][3][2] , \s_mX2[0][3][1] , 
        \s_mX2[0][3][0] }) );
  Mux_NBit_2x1_NBIT_IN8_4 MUX4_3_1 ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .port1({n9, n12, s_msb[5:3], n7, n15, n8}), .sel(
        n21), .portY({\s_mX2[0][3][15] , \s_mX2[0][3][14] , \s_mX2[0][3][13] , 
        \s_mX2[0][3][12] , \s_mX2[0][3][11] , \s_mX2[0][3][10] , 
        \s_mX2[0][3][9] , \s_mX2[0][3][8] }) );
  Mux_NBit_2x1_NBIT_IN8_3 MUX4_3_2 ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .port1({s_msb[7:3], n7, s_msb[1], n8}), .sel(n20), 
        .portY({\s_mX2[0][3][23] , \s_mX2[0][3][22] , \s_mX2[0][3][21] , 
        \s_mX2[0][3][20] , \s_mX2[0][3][19] , \s_mX2[0][3][18] , 
        \s_mX2[0][3][17] , \s_mX2[0][3][16] }) );
  Mux_NBit_2x1_NBIT_IN8_2 MUX4_3_3 ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .port1(s_msb), .sel(n20), .portY({
        \s_mX2[0][3][31] , \s_mX2[0][3][30] , \s_mX2[0][3][29] , 
        \s_mX2[0][3][28] , \s_mX2[0][3][27] , \s_mX2[0][3][26] , 
        \s_mX2[0][3][25] , \s_mX2[0][3][24] }) );
  Mux_NBit_2x1_NBIT_IN8_1 MUX3_3_4 ( .port0(BS_data_in[7:0]), .port1(s_msb), 
        .sel(n20), .portY({\s_mX2[0][3][39] , \s_mX2[0][3][38] , 
        \s_mX2[0][3][37] , \s_mX2[0][3][36] , \s_mX2[0][3][35] , 
        \s_mX2[0][3][34] , \s_mX2[0][3][33] , \s_mX2[0][3][32] }) );
  Mux_NBit_2x1_NBIT_IN40_0 MUX1_0_0 ( .port0({\s_mX2[0][0][39] , 
        \s_mX2[0][0][38] , \s_mX2[0][0][37] , \s_mX2[0][0][36] , 
        \s_mX2[0][0][35] , \s_mX2[0][0][34] , \s_mX2[0][0][33] , 
        \s_mX2[0][0][32] , \s_mX2[0][0][31] , \s_mX2[0][0][30] , 
        \s_mX2[0][0][29] , \s_mX2[0][0][28] , \s_mX2[0][0][27] , 
        \s_mX2[0][0][26] , \s_mX2[0][0][25] , \s_mX2[0][0][24] , 
        \s_mX2[0][0][23] , \s_mX2[0][0][22] , \s_mX2[0][0][21] , 
        \s_mX2[0][0][20] , \s_mX2[0][0][19] , \s_mX2[0][0][18] , 
        \s_mX2[0][0][17] , \s_mX2[0][0][16] , \s_mX2[0][0][15] , 
        \s_mX2[0][0][14] , \s_mX2[0][0][13] , \s_mX2[0][0][12] , 
        \s_mX2[0][0][11] , \s_mX2[0][0][10] , \s_mX2[0][0][9] , 
        \s_mX2[0][0][8] , \s_mX2[0][0][7] , \s_mX2[0][0][6] , \s_mX2[0][0][5] , 
        \s_mX2[0][0][4] , \s_mX2[0][0][3] , \s_mX2[0][0][2] , \s_mX2[0][0][1] , 
        \s_mX2[0][0][0] }), .port1({\s_mX2[0][1][39] , \s_mX2[0][1][38] , 
        \s_mX2[0][1][37] , \s_mX2[0][1][36] , \s_mX2[0][1][35] , 
        \s_mX2[0][1][34] , \s_mX2[0][1][33] , \s_mX2[0][1][32] , 
        \s_mX2[0][1][31] , \s_mX2[0][1][30] , \s_mX2[0][1][29] , 
        \s_mX2[0][1][28] , \s_mX2[0][1][27] , \s_mX2[0][1][26] , 
        \s_mX2[0][1][25] , \s_mX2[0][1][24] , \s_mX2[0][1][23] , 
        \s_mX2[0][1][22] , \s_mX2[0][1][21] , \s_mX2[0][1][20] , 
        \s_mX2[0][1][19] , \s_mX2[0][1][18] , \s_mX2[0][1][17] , 
        \s_mX2[0][1][16] , \s_mX2[0][1][15] , \s_mX2[0][1][14] , 
        \s_mX2[0][1][13] , \s_mX2[0][1][12] , \s_mX2[0][1][11] , 
        \s_mX2[0][1][10] , \s_mX2[0][1][9] , \s_mX2[0][1][8] , 
        \s_mX2[0][1][7] , \s_mX2[0][1][6] , \s_mX2[0][1][5] , \s_mX2[0][1][4] , 
        \s_mX2[0][1][3] , \s_mX2[0][1][2] , \s_mX2[0][1][1] , \s_mX2[0][1][0] }), .sel(BS_amount[3]), .portY({\s_mX2[1][0][39] , \s_mX2[1][0][38] , 
        \s_mX2[1][0][37] , \s_mX2[1][0][36] , \s_mX2[1][0][35] , 
        \s_mX2[1][0][34] , \s_mX2[1][0][33] , \s_mX2[1][0][32] , 
        \s_mX2[1][0][31] , \s_mX2[1][0][30] , \s_mX2[1][0][29] , 
        \s_mX2[1][0][28] , \s_mX2[1][0][27] , \s_mX2[1][0][26] , 
        \s_mX2[1][0][25] , \s_mX2[1][0][24] , \s_mX2[1][0][23] , 
        \s_mX2[1][0][22] , \s_mX2[1][0][21] , \s_mX2[1][0][20] , 
        \s_mX2[1][0][19] , \s_mX2[1][0][18] , \s_mX2[1][0][17] , 
        \s_mX2[1][0][16] , \s_mX2[1][0][15] , \s_mX2[1][0][14] , 
        \s_mX2[1][0][13] , \s_mX2[1][0][12] , \s_mX2[1][0][11] , 
        \s_mX2[1][0][10] , \s_mX2[1][0][9] , \s_mX2[1][0][8] , 
        \s_mX2[1][0][7] , \s_mX2[1][0][6] , \s_mX2[1][0][5] , \s_mX2[1][0][4] , 
        \s_mX2[1][0][3] , \s_mX2[1][0][2] , \s_mX2[1][0][1] , \s_mX2[1][0][0] }) );
  Mux_NBit_2x1_NBIT_IN40_3 MUX1_0_2_0 ( .port0({\s_mX2[0][2][39] , 
        \s_mX2[0][2][38] , \s_mX2[0][2][37] , \s_mX2[0][2][36] , 
        \s_mX2[0][2][35] , \s_mX2[0][2][34] , \s_mX2[0][2][33] , 
        \s_mX2[0][2][32] , \s_mX2[0][2][31] , \s_mX2[0][2][30] , 
        \s_mX2[0][2][29] , \s_mX2[0][2][28] , \s_mX2[0][2][27] , 
        \s_mX2[0][2][26] , \s_mX2[0][2][25] , \s_mX2[0][2][24] , 
        \s_mX2[0][2][23] , \s_mX2[0][2][22] , \s_mX2[0][2][21] , 
        \s_mX2[0][2][20] , \s_mX2[0][2][19] , \s_mX2[0][2][18] , 
        \s_mX2[0][2][17] , \s_mX2[0][2][16] , \s_mX2[0][2][15] , 
        \s_mX2[0][2][14] , \s_mX2[0][2][13] , \s_mX2[0][2][12] , 
        \s_mX2[0][2][11] , \s_mX2[0][2][10] , \s_mX2[0][2][9] , 
        \s_mX2[0][2][8] , \s_mX2[0][2][7] , \s_mX2[0][2][6] , \s_mX2[0][2][5] , 
        \s_mX2[0][2][4] , \s_mX2[0][2][3] , \s_mX2[0][2][2] , \s_mX2[0][2][1] , 
        \s_mX2[0][2][0] }), .port1({\s_mX2[0][3][39] , \s_mX2[0][3][38] , 
        \s_mX2[0][3][37] , \s_mX2[0][3][36] , \s_mX2[0][3][35] , 
        \s_mX2[0][3][34] , \s_mX2[0][3][33] , \s_mX2[0][3][32] , 
        \s_mX2[0][3][31] , \s_mX2[0][3][30] , \s_mX2[0][3][29] , 
        \s_mX2[0][3][28] , \s_mX2[0][3][27] , \s_mX2[0][3][26] , 
        \s_mX2[0][3][25] , \s_mX2[0][3][24] , \s_mX2[0][3][23] , 
        \s_mX2[0][3][22] , \s_mX2[0][3][21] , \s_mX2[0][3][20] , 
        \s_mX2[0][3][19] , \s_mX2[0][3][18] , \s_mX2[0][3][17] , 
        \s_mX2[0][3][16] , \s_mX2[0][3][15] , \s_mX2[0][3][14] , 
        \s_mX2[0][3][13] , \s_mX2[0][3][12] , \s_mX2[0][3][11] , 
        \s_mX2[0][3][10] , \s_mX2[0][3][9] , \s_mX2[0][3][8] , 
        \s_mX2[0][3][7] , \s_mX2[0][3][6] , \s_mX2[0][3][5] , \s_mX2[0][3][4] , 
        \s_mX2[0][3][3] , \s_mX2[0][3][2] , \s_mX2[0][3][1] , \s_mX2[0][3][0] }), .sel(BS_amount[3]), .portY({\s_mX2[1][2][39] , \s_mX2[1][2][38] , 
        \s_mX2[1][2][37] , \s_mX2[1][2][36] , \s_mX2[1][2][35] , 
        \s_mX2[1][2][34] , \s_mX2[1][2][33] , \s_mX2[1][2][32] , 
        \s_mX2[1][2][31] , \s_mX2[1][2][30] , \s_mX2[1][2][29] , 
        \s_mX2[1][2][28] , \s_mX2[1][2][27] , \s_mX2[1][2][26] , 
        \s_mX2[1][2][25] , \s_mX2[1][2][24] , \s_mX2[1][2][23] , 
        \s_mX2[1][2][22] , \s_mX2[1][2][21] , \s_mX2[1][2][20] , 
        \s_mX2[1][2][19] , \s_mX2[1][2][18] , \s_mX2[1][2][17] , 
        \s_mX2[1][2][16] , \s_mX2[1][2][15] , \s_mX2[1][2][14] , 
        \s_mX2[1][2][13] , \s_mX2[1][2][12] , \s_mX2[1][2][11] , 
        \s_mX2[1][2][10] , \s_mX2[1][2][9] , \s_mX2[1][2][8] , 
        \s_mX2[1][2][7] , \s_mX2[1][2][6] , \s_mX2[1][2][5] , \s_mX2[1][2][4] , 
        \s_mX2[1][2][3] , \s_mX2[1][2][2] , \s_mX2[1][2][1] , \s_mX2[1][2][0] }) );
  Mux_NBit_2x1_NBIT_IN40_2 MUX1_1_0 ( .port0({\s_mX2[1][0][39] , 
        \s_mX2[1][0][38] , \s_mX2[1][0][37] , \s_mX2[1][0][36] , 
        \s_mX2[1][0][35] , \s_mX2[1][0][34] , \s_mX2[1][0][33] , 
        \s_mX2[1][0][32] , \s_mX2[1][0][31] , \s_mX2[1][0][30] , 
        \s_mX2[1][0][29] , \s_mX2[1][0][28] , \s_mX2[1][0][27] , 
        \s_mX2[1][0][26] , \s_mX2[1][0][25] , \s_mX2[1][0][24] , 
        \s_mX2[1][0][23] , \s_mX2[1][0][22] , \s_mX2[1][0][21] , 
        \s_mX2[1][0][20] , \s_mX2[1][0][19] , \s_mX2[1][0][18] , 
        \s_mX2[1][0][17] , \s_mX2[1][0][16] , \s_mX2[1][0][15] , 
        \s_mX2[1][0][14] , \s_mX2[1][0][13] , \s_mX2[1][0][12] , 
        \s_mX2[1][0][11] , \s_mX2[1][0][10] , \s_mX2[1][0][9] , 
        \s_mX2[1][0][8] , \s_mX2[1][0][7] , \s_mX2[1][0][6] , \s_mX2[1][0][5] , 
        \s_mX2[1][0][4] , \s_mX2[1][0][3] , \s_mX2[1][0][2] , \s_mX2[1][0][1] , 
        \s_mX2[1][0][0] }), .port1({\s_mX2[1][2][39] , \s_mX2[1][2][38] , 
        \s_mX2[1][2][37] , \s_mX2[1][2][36] , \s_mX2[1][2][35] , 
        \s_mX2[1][2][34] , \s_mX2[1][2][33] , \s_mX2[1][2][32] , 
        \s_mX2[1][2][31] , \s_mX2[1][2][30] , \s_mX2[1][2][29] , 
        \s_mX2[1][2][28] , \s_mX2[1][2][27] , \s_mX2[1][2][26] , 
        \s_mX2[1][2][25] , \s_mX2[1][2][24] , \s_mX2[1][2][23] , 
        \s_mX2[1][2][22] , \s_mX2[1][2][21] , \s_mX2[1][2][20] , 
        \s_mX2[1][2][19] , \s_mX2[1][2][18] , \s_mX2[1][2][17] , 
        \s_mX2[1][2][16] , \s_mX2[1][2][15] , \s_mX2[1][2][14] , 
        \s_mX2[1][2][13] , \s_mX2[1][2][12] , \s_mX2[1][2][11] , 
        \s_mX2[1][2][10] , \s_mX2[1][2][9] , \s_mX2[1][2][8] , 
        \s_mX2[1][2][7] , \s_mX2[1][2][6] , \s_mX2[1][2][5] , \s_mX2[1][2][4] , 
        \s_mX2[1][2][3] , \s_mX2[1][2][2] , \s_mX2[1][2][1] , \s_mX2[1][2][0] }), .sel(BS_amount[4]), .portY({\s_mX2[2][0][39] , \s_mX2[2][0][38] , 
        \s_mX2[2][0][37] , \s_mX2[2][0][36] , \s_mX2[2][0][35] , 
        \s_mX2[2][0][34] , \s_mX2[2][0][33] , \s_mX2[2][0][32] , 
        \s_mX2[2][0][31] , \s_mX2[2][0][30] , \s_mX2[2][0][29] , 
        \s_mX2[2][0][28] , \s_mX2[2][0][27] , \s_mX2[2][0][26] , 
        \s_mX2[2][0][25] , \s_mX2[2][0][24] , \s_mX2[2][0][23] , 
        \s_mX2[2][0][22] , \s_mX2[2][0][21] , \s_mX2[2][0][20] , 
        \s_mX2[2][0][19] , \s_mX2[2][0][18] , \s_mX2[2][0][17] , 
        \s_mX2[2][0][16] , \s_mX2[2][0][15] , \s_mX2[2][0][14] , 
        \s_mX2[2][0][13] , \s_mX2[2][0][12] , \s_mX2[2][0][11] , 
        \s_mX2[2][0][10] , \s_mX2[2][0][9] , \s_mX2[2][0][8] , 
        \s_mX2[2][0][7] , \s_mX2[2][0][6] , \s_mX2[2][0][5] , \s_mX2[2][0][4] , 
        \s_mX2[2][0][3] , \s_mX2[2][0][2] , \s_mX2[2][0][1] , \s_mX2[2][0][0] }) );
  Mux_NBit_2x1_NBIT_IN40_1 MUX_selected_mask ( .port0({\s_mX2[2][0][39] , 
        \s_mX2[2][0][38] , \s_mX2[2][0][37] , \s_mX2[2][0][36] , 
        \s_mX2[2][0][35] , \s_mX2[2][0][34] , \s_mX2[2][0][33] , 
        \s_mX2[2][0][32] , \s_mX2[2][0][31] , n13, \s_mX2[2][0][29] , 
        \s_mX2[2][0][28] , \s_mX2[2][0][27] , \s_mX2[2][0][26] , 
        \s_mX2[2][0][25] , \s_mX2[2][0][24] , \s_mX2[2][0][23] , 
        \s_mX2[2][0][22] , \s_mX2[2][0][21] , \s_mX2[2][0][20] , 
        \s_mX2[2][0][19] , \s_mX2[2][0][18] , \s_mX2[2][0][17] , 
        \s_mX2[2][0][16] , \s_mX2[2][0][15] , \s_mX2[2][0][14] , 
        \s_mX2[2][0][13] , \s_mX2[2][0][12] , \s_mX2[2][0][11] , 
        \s_mX2[2][0][10] , \s_mX2[2][0][9] , \s_mX2[2][0][8] , 
        \s_mX2[2][0][7] , \s_mX2[2][0][6] , \s_mX2[2][0][5] , \s_mX2[2][0][4] , 
        \s_mX2[2][0][3] , \s_mX2[2][0][2] , \s_mX2[2][0][1] , \s_mX2[2][0][0] }), .port1({\s_mX2[2][0][38] , \s_mX2[2][0][37] , \s_mX2[2][0][36] , 
        \s_mX2[2][0][35] , \s_mX2[2][0][34] , \s_mX2[2][0][33] , 
        \s_mX2[2][0][32] , \s_mX2[2][0][31] , \s_mX2[2][0][30] , 
        \s_mX2[2][0][29] , \s_mX2[2][0][28] , \s_mX2[2][0][27] , 
        \s_mX2[2][0][26] , \s_mX2[2][0][25] , \s_mX2[2][0][24] , 
        \s_mX2[2][0][23] , \s_mX2[2][0][22] , \s_mX2[2][0][21] , 
        \s_mX2[2][0][20] , \s_mX2[2][0][19] , \s_mX2[2][0][18] , 
        \s_mX2[2][0][17] , \s_mX2[2][0][16] , \s_mX2[2][0][15] , 
        \s_mX2[2][0][14] , \s_mX2[2][0][13] , \s_mX2[2][0][12] , 
        \s_mX2[2][0][11] , \s_mX2[2][0][10] , \s_mX2[2][0][9] , 
        \s_mX2[2][0][8] , \s_mX2[2][0][7] , \s_mX2[2][0][6] , \s_mX2[2][0][5] , 
        \s_mX2[2][0][4] , \s_mX2[2][0][3] , \s_mX2[2][0][2] , \s_mX2[2][0][1] , 
        \s_mX2[2][0][0] , 1'b0}), .sel(n26), .portY({s_selected_mask, 
        SYNOPSYS_UNCONNECTED__0}) );
  Mux_NBit_2x1_NBIT_IN3 MUX3x1 ( .port0(s_amount), .port1(s_not_amount), .sel(
        n26), .portY(s_sel_out) );
  Mux_NBit_2x1_NBIT_IN32_7 MUX2_0_0_0 ( .port0({s_selected_mask[39:35], n14, 
        s_selected_mask[33], n16, n11, s_selected_mask[30:8]}), .port1({
        s_selected_mask[38:33], n16, n11, s_selected_mask[30:7]}), .sel(
        s_sel_out[0]), .portY({\s_out_mask[1][0][31] , \s_out_mask[1][0][30] , 
        \s_out_mask[1][0][29] , \s_out_mask[1][0][28] , \s_out_mask[1][0][27] , 
        \s_out_mask[1][0][26] , \s_out_mask[1][0][25] , \s_out_mask[1][0][24] , 
        \s_out_mask[1][0][23] , \s_out_mask[1][0][22] , \s_out_mask[1][0][21] , 
        \s_out_mask[1][0][20] , \s_out_mask[1][0][19] , \s_out_mask[1][0][18] , 
        \s_out_mask[1][0][17] , \s_out_mask[1][0][16] , \s_out_mask[1][0][15] , 
        \s_out_mask[1][0][14] , \s_out_mask[1][0][13] , \s_out_mask[1][0][12] , 
        \s_out_mask[1][0][11] , \s_out_mask[1][0][10] , \s_out_mask[1][0][9] , 
        \s_out_mask[1][0][8] , \s_out_mask[1][0][7] , \s_out_mask[1][0][6] , 
        \s_out_mask[1][0][5] , \s_out_mask[1][0][4] , \s_out_mask[1][0][3] , 
        \s_out_mask[1][0][2] , \s_out_mask[1][0][1] , \s_out_mask[1][0][0] })
         );
  Mux_NBit_2x1_NBIT_IN32_6 MUX2_0_2 ( .port0({s_selected_mask[37:33], n16, n11, 
        s_selected_mask[30:6]}), .port1({s_selected_mask[36:32], n6, 
        s_selected_mask[30:5]}), .sel(s_sel_out[0]), .portY({
        \s_out_mask[1][2][31] , \s_out_mask[1][2][30] , \s_out_mask[1][2][29] , 
        \s_out_mask[1][2][28] , \s_out_mask[1][2][27] , \s_out_mask[1][2][26] , 
        \s_out_mask[1][2][25] , \s_out_mask[1][2][24] , \s_out_mask[1][2][23] , 
        \s_out_mask[1][2][22] , \s_out_mask[1][2][21] , \s_out_mask[1][2][20] , 
        \s_out_mask[1][2][19] , \s_out_mask[1][2][18] , \s_out_mask[1][2][17] , 
        \s_out_mask[1][2][16] , \s_out_mask[1][2][15] , \s_out_mask[1][2][14] , 
        \s_out_mask[1][2][13] , \s_out_mask[1][2][12] , \s_out_mask[1][2][11] , 
        \s_out_mask[1][2][10] , \s_out_mask[1][2][9] , \s_out_mask[1][2][8] , 
        \s_out_mask[1][2][7] , \s_out_mask[1][2][6] , \s_out_mask[1][2][5] , 
        \s_out_mask[1][2][4] , \s_out_mask[1][2][3] , \s_out_mask[1][2][2] , 
        \s_out_mask[1][2][1] , \s_out_mask[1][2][0] }) );
  Mux_NBit_2x1_NBIT_IN32_5 MUX2_0_4 ( .port0(s_selected_mask[35:4]), .port1(
        s_selected_mask[34:3]), .sel(s_sel_out[0]), .portY({
        \s_out_mask[1][4][31] , \s_out_mask[1][4][30] , \s_out_mask[1][4][29] , 
        \s_out_mask[1][4][28] , \s_out_mask[1][4][27] , \s_out_mask[1][4][26] , 
        \s_out_mask[1][4][25] , \s_out_mask[1][4][24] , \s_out_mask[1][4][23] , 
        \s_out_mask[1][4][22] , \s_out_mask[1][4][21] , \s_out_mask[1][4][20] , 
        \s_out_mask[1][4][19] , \s_out_mask[1][4][18] , \s_out_mask[1][4][17] , 
        \s_out_mask[1][4][16] , \s_out_mask[1][4][15] , \s_out_mask[1][4][14] , 
        \s_out_mask[1][4][13] , \s_out_mask[1][4][12] , \s_out_mask[1][4][11] , 
        \s_out_mask[1][4][10] , \s_out_mask[1][4][9] , \s_out_mask[1][4][8] , 
        \s_out_mask[1][4][7] , \s_out_mask[1][4][6] , \s_out_mask[1][4][5] , 
        \s_out_mask[1][4][4] , \s_out_mask[1][4][3] , \s_out_mask[1][4][2] , 
        \s_out_mask[1][4][1] , \s_out_mask[1][4][0] }) );
  Mux_NBit_2x1_NBIT_IN32_4 MUX2_0_6 ( .port0(s_selected_mask[33:2]), .port1(
        s_selected_mask[32:1]), .sel(s_sel_out[0]), .portY({
        \s_out_mask[1][6][31] , \s_out_mask[1][6][30] , \s_out_mask[1][6][29] , 
        \s_out_mask[1][6][28] , \s_out_mask[1][6][27] , \s_out_mask[1][6][26] , 
        \s_out_mask[1][6][25] , \s_out_mask[1][6][24] , \s_out_mask[1][6][23] , 
        \s_out_mask[1][6][22] , \s_out_mask[1][6][21] , \s_out_mask[1][6][20] , 
        \s_out_mask[1][6][19] , \s_out_mask[1][6][18] , \s_out_mask[1][6][17] , 
        \s_out_mask[1][6][16] , \s_out_mask[1][6][15] , \s_out_mask[1][6][14] , 
        \s_out_mask[1][6][13] , \s_out_mask[1][6][12] , \s_out_mask[1][6][11] , 
        \s_out_mask[1][6][10] , \s_out_mask[1][6][9] , \s_out_mask[1][6][8] , 
        \s_out_mask[1][6][7] , \s_out_mask[1][6][6] , \s_out_mask[1][6][5] , 
        \s_out_mask[1][6][4] , \s_out_mask[1][6][3] , \s_out_mask[1][6][2] , 
        \s_out_mask[1][6][1] , \s_out_mask[1][6][0] }) );
  Mux_NBit_2x1_NBIT_IN32_3 MUX2_1_0_0 ( .port0({\s_out_mask[1][0][31] , 
        \s_out_mask[1][0][30] , \s_out_mask[1][0][29] , \s_out_mask[1][0][28] , 
        \s_out_mask[1][0][27] , \s_out_mask[1][0][26] , \s_out_mask[1][0][25] , 
        \s_out_mask[1][0][24] , \s_out_mask[1][0][23] , \s_out_mask[1][0][22] , 
        \s_out_mask[1][0][21] , \s_out_mask[1][0][20] , \s_out_mask[1][0][19] , 
        \s_out_mask[1][0][18] , \s_out_mask[1][0][17] , \s_out_mask[1][0][16] , 
        \s_out_mask[1][0][15] , \s_out_mask[1][0][14] , \s_out_mask[1][0][13] , 
        \s_out_mask[1][0][12] , \s_out_mask[1][0][11] , \s_out_mask[1][0][10] , 
        \s_out_mask[1][0][9] , \s_out_mask[1][0][8] , \s_out_mask[1][0][7] , 
        \s_out_mask[1][0][6] , \s_out_mask[1][0][5] , \s_out_mask[1][0][4] , 
        \s_out_mask[1][0][3] , \s_out_mask[1][0][2] , \s_out_mask[1][0][1] , 
        \s_out_mask[1][0][0] }), .port1({\s_out_mask[1][2][31] , 
        \s_out_mask[1][2][30] , \s_out_mask[1][2][29] , \s_out_mask[1][2][28] , 
        \s_out_mask[1][2][27] , \s_out_mask[1][2][26] , \s_out_mask[1][2][25] , 
        \s_out_mask[1][2][24] , \s_out_mask[1][2][23] , \s_out_mask[1][2][22] , 
        \s_out_mask[1][2][21] , \s_out_mask[1][2][20] , \s_out_mask[1][2][19] , 
        \s_out_mask[1][2][18] , \s_out_mask[1][2][17] , \s_out_mask[1][2][16] , 
        \s_out_mask[1][2][15] , \s_out_mask[1][2][14] , \s_out_mask[1][2][13] , 
        \s_out_mask[1][2][12] , \s_out_mask[1][2][11] , \s_out_mask[1][2][10] , 
        \s_out_mask[1][2][9] , \s_out_mask[1][2][8] , \s_out_mask[1][2][7] , 
        \s_out_mask[1][2][6] , \s_out_mask[1][2][5] , \s_out_mask[1][2][4] , 
        \s_out_mask[1][2][3] , \s_out_mask[1][2][2] , \s_out_mask[1][2][1] , 
        \s_out_mask[1][2][0] }), .sel(s_sel_out[1]), .portY({
        \s_out_mask[2][0][31] , \s_out_mask[2][0][30] , \s_out_mask[2][0][29] , 
        \s_out_mask[2][0][28] , \s_out_mask[2][0][27] , \s_out_mask[2][0][26] , 
        \s_out_mask[2][0][25] , \s_out_mask[2][0][24] , \s_out_mask[2][0][23] , 
        \s_out_mask[2][0][22] , \s_out_mask[2][0][21] , \s_out_mask[2][0][20] , 
        \s_out_mask[2][0][19] , \s_out_mask[2][0][18] , \s_out_mask[2][0][17] , 
        \s_out_mask[2][0][16] , \s_out_mask[2][0][15] , \s_out_mask[2][0][14] , 
        \s_out_mask[2][0][13] , \s_out_mask[2][0][12] , \s_out_mask[2][0][11] , 
        \s_out_mask[2][0][10] , \s_out_mask[2][0][9] , \s_out_mask[2][0][8] , 
        \s_out_mask[2][0][7] , \s_out_mask[2][0][6] , \s_out_mask[2][0][5] , 
        \s_out_mask[2][0][4] , \s_out_mask[2][0][3] , \s_out_mask[2][0][2] , 
        \s_out_mask[2][0][1] , \s_out_mask[2][0][0] }) );
  Mux_NBit_2x1_NBIT_IN32_2 MUX2_1_4 ( .port0({\s_out_mask[1][4][31] , 
        \s_out_mask[1][4][30] , \s_out_mask[1][4][29] , \s_out_mask[1][4][28] , 
        \s_out_mask[1][4][27] , \s_out_mask[1][4][26] , \s_out_mask[1][4][25] , 
        \s_out_mask[1][4][24] , \s_out_mask[1][4][23] , \s_out_mask[1][4][22] , 
        \s_out_mask[1][4][21] , \s_out_mask[1][4][20] , \s_out_mask[1][4][19] , 
        \s_out_mask[1][4][18] , \s_out_mask[1][4][17] , \s_out_mask[1][4][16] , 
        \s_out_mask[1][4][15] , \s_out_mask[1][4][14] , \s_out_mask[1][4][13] , 
        \s_out_mask[1][4][12] , \s_out_mask[1][4][11] , \s_out_mask[1][4][10] , 
        \s_out_mask[1][4][9] , \s_out_mask[1][4][8] , \s_out_mask[1][4][7] , 
        \s_out_mask[1][4][6] , \s_out_mask[1][4][5] , \s_out_mask[1][4][4] , 
        \s_out_mask[1][4][3] , \s_out_mask[1][4][2] , \s_out_mask[1][4][1] , 
        \s_out_mask[1][4][0] }), .port1({\s_out_mask[1][6][31] , 
        \s_out_mask[1][6][30] , \s_out_mask[1][6][29] , \s_out_mask[1][6][28] , 
        \s_out_mask[1][6][27] , \s_out_mask[1][6][26] , \s_out_mask[1][6][25] , 
        \s_out_mask[1][6][24] , \s_out_mask[1][6][23] , \s_out_mask[1][6][22] , 
        \s_out_mask[1][6][21] , \s_out_mask[1][6][20] , \s_out_mask[1][6][19] , 
        \s_out_mask[1][6][18] , \s_out_mask[1][6][17] , \s_out_mask[1][6][16] , 
        \s_out_mask[1][6][15] , \s_out_mask[1][6][14] , \s_out_mask[1][6][13] , 
        \s_out_mask[1][6][12] , \s_out_mask[1][6][11] , \s_out_mask[1][6][10] , 
        \s_out_mask[1][6][9] , \s_out_mask[1][6][8] , \s_out_mask[1][6][7] , 
        \s_out_mask[1][6][6] , \s_out_mask[1][6][5] , \s_out_mask[1][6][4] , 
        \s_out_mask[1][6][3] , \s_out_mask[1][6][2] , \s_out_mask[1][6][1] , 
        \s_out_mask[1][6][0] }), .sel(s_sel_out[1]), .portY({
        \s_out_mask[2][4][31] , \s_out_mask[2][4][30] , \s_out_mask[2][4][29] , 
        \s_out_mask[2][4][28] , \s_out_mask[2][4][27] , \s_out_mask[2][4][26] , 
        \s_out_mask[2][4][25] , \s_out_mask[2][4][24] , \s_out_mask[2][4][23] , 
        \s_out_mask[2][4][22] , \s_out_mask[2][4][21] , \s_out_mask[2][4][20] , 
        \s_out_mask[2][4][19] , \s_out_mask[2][4][18] , \s_out_mask[2][4][17] , 
        \s_out_mask[2][4][16] , \s_out_mask[2][4][15] , \s_out_mask[2][4][14] , 
        \s_out_mask[2][4][13] , \s_out_mask[2][4][12] , \s_out_mask[2][4][11] , 
        \s_out_mask[2][4][10] , \s_out_mask[2][4][9] , \s_out_mask[2][4][8] , 
        \s_out_mask[2][4][7] , \s_out_mask[2][4][6] , \s_out_mask[2][4][5] , 
        \s_out_mask[2][4][4] , \s_out_mask[2][4][3] , \s_out_mask[2][4][2] , 
        \s_out_mask[2][4][1] , \s_out_mask[2][4][0] }) );
  Mux_NBit_2x1_NBIT_IN32_1 MUX2_2_0_0 ( .port0({\s_out_mask[2][0][31] , 
        \s_out_mask[2][0][30] , \s_out_mask[2][0][29] , \s_out_mask[2][0][28] , 
        \s_out_mask[2][0][27] , \s_out_mask[2][0][26] , \s_out_mask[2][0][25] , 
        \s_out_mask[2][0][24] , \s_out_mask[2][0][23] , \s_out_mask[2][0][22] , 
        \s_out_mask[2][0][21] , \s_out_mask[2][0][20] , \s_out_mask[2][0][19] , 
        \s_out_mask[2][0][18] , \s_out_mask[2][0][17] , \s_out_mask[2][0][16] , 
        \s_out_mask[2][0][15] , \s_out_mask[2][0][14] , \s_out_mask[2][0][13] , 
        \s_out_mask[2][0][12] , \s_out_mask[2][0][11] , \s_out_mask[2][0][10] , 
        \s_out_mask[2][0][9] , \s_out_mask[2][0][8] , \s_out_mask[2][0][7] , 
        \s_out_mask[2][0][6] , \s_out_mask[2][0][5] , \s_out_mask[2][0][4] , 
        \s_out_mask[2][0][3] , \s_out_mask[2][0][2] , \s_out_mask[2][0][1] , 
        \s_out_mask[2][0][0] }), .port1({\s_out_mask[2][4][31] , 
        \s_out_mask[2][4][30] , \s_out_mask[2][4][29] , \s_out_mask[2][4][28] , 
        \s_out_mask[2][4][27] , \s_out_mask[2][4][26] , \s_out_mask[2][4][25] , 
        \s_out_mask[2][4][24] , \s_out_mask[2][4][23] , \s_out_mask[2][4][22] , 
        \s_out_mask[2][4][21] , \s_out_mask[2][4][20] , \s_out_mask[2][4][19] , 
        \s_out_mask[2][4][18] , \s_out_mask[2][4][17] , \s_out_mask[2][4][16] , 
        \s_out_mask[2][4][15] , \s_out_mask[2][4][14] , \s_out_mask[2][4][13] , 
        \s_out_mask[2][4][12] , \s_out_mask[2][4][11] , \s_out_mask[2][4][10] , 
        \s_out_mask[2][4][9] , \s_out_mask[2][4][8] , \s_out_mask[2][4][7] , 
        \s_out_mask[2][4][6] , \s_out_mask[2][4][5] , \s_out_mask[2][4][4] , 
        \s_out_mask[2][4][3] , \s_out_mask[2][4][2] , \s_out_mask[2][4][1] , 
        \s_out_mask[2][4][0] }), .sel(s_sel_out[2]), .portY(BS_data_out) );
  CLKBUF_X1 U2 ( .A(s_selected_mask[31]), .Z(n6) );
  CLKBUF_X1 U3 ( .A(s_msb[2]), .Z(n7) );
  CLKBUF_X1 U4 ( .A(s_msb[0]), .Z(n8) );
  CLKBUF_X1 U5 ( .A(s_msb[7]), .Z(n9) );
  CLKBUF_X1 U6 ( .A(BS_data_in[31]), .Z(n10) );
  CLKBUF_X1 U7 ( .A(n6), .Z(n11) );
  CLKBUF_X1 U8 ( .A(s_msb[6]), .Z(n12) );
  BUF_X2 U9 ( .A(n18), .Z(n25) );
  BUF_X2 U10 ( .A(n18), .Z(n24) );
  BUF_X2 U11 ( .A(n17), .Z(n22) );
  BUF_X2 U12 ( .A(n17), .Z(n20) );
  BUF_X1 U13 ( .A(n17), .Z(n21) );
  BUF_X1 U14 ( .A(n18), .Z(n23) );
  OR2_X1 U15 ( .A1(BS_opcode[1]), .A2(n19), .ZN(n5) );
  BUF_X1 U16 ( .A(n4), .Z(n18) );
  BUF_X1 U17 ( .A(n4), .Z(n17) );
  CLKBUF_X1 U18 ( .A(n4), .Z(n19) );
  INV_X1 U19 ( .A(s_not_amount[0]), .ZN(s_amount[0]) );
  INV_X1 U20 ( .A(s_not_amount[1]), .ZN(s_amount[1]) );
  NAND2_X1 U21 ( .A1(BS_amount[1]), .A2(n5), .ZN(s_not_amount[1]) );
  INV_X1 U22 ( .A(s_not_amount[2]), .ZN(s_amount[2]) );
  NAND2_X1 U23 ( .A1(BS_amount[2]), .A2(n5), .ZN(s_not_amount[2]) );
  CLKBUF_X1 U24 ( .A(\s_mX2[2][0][30] ), .Z(n13) );
  CLKBUF_X1 U25 ( .A(s_selected_mask[34]), .Z(n14) );
  CLKBUF_X1 U26 ( .A(s_msb[1]), .Z(n15) );
  CLKBUF_X1 U27 ( .A(s_selected_mask[32]), .Z(n16) );
  NAND2_X1 U28 ( .A1(BS_amount[0]), .A2(n5), .ZN(s_not_amount[0]) );
  CLKBUF_X3 U29 ( .A(n19), .Z(n26) );
endmodule


module Mux_NBit_2x1_NBIT_IN6_0 ( port0, port1, sel, portY );
  input [5:0] port0;
  input [5:0] port1;
  output [5:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, n8, n9, n10, n11, n12, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;

  INV_X1 U1 ( .A(sel), .ZN(n9) );
  INV_X1 U2 ( .A(n8), .ZN(N7) );
  AOI22_X1 U3 ( .A1(port0[5]), .A2(n9), .B1(sel), .B2(port1[5]), .ZN(n8) );
  INV_X1 U4 ( .A(n14), .ZN(N2) );
  AOI22_X1 U5 ( .A1(port0[0]), .A2(n9), .B1(port1[0]), .B2(sel), .ZN(n14) );
  INV_X1 U6 ( .A(n13), .ZN(N3) );
  AOI22_X1 U7 ( .A1(port0[1]), .A2(n9), .B1(port1[1]), .B2(sel), .ZN(n13) );
  INV_X1 U8 ( .A(n12), .ZN(N4) );
  AOI22_X1 U9 ( .A1(port0[2]), .A2(n9), .B1(port1[2]), .B2(sel), .ZN(n12) );
  INV_X1 U10 ( .A(n11), .ZN(N5) );
  AOI22_X1 U11 ( .A1(port0[3]), .A2(n9), .B1(port1[3]), .B2(sel), .ZN(n11) );
  INV_X1 U12 ( .A(n10), .ZN(N6) );
  AOI22_X1 U13 ( .A1(port0[4]), .A2(n9), .B1(port1[4]), .B2(sel), .ZN(n10) );
endmodule


module Mux_NBit_2x1_NBIT_IN10_0 ( port0, port1, sel, portY );
  input [9:0] port0;
  input [9:0] port1;
  output [9:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;

  INV_X1 U1 ( .A(sel), .ZN(n13) );
  INV_X1 U2 ( .A(n16), .ZN(N6) );
  AOI22_X1 U3 ( .A1(port0[4]), .A2(n13), .B1(port1[4]), .B2(sel), .ZN(n16) );
  INV_X1 U4 ( .A(n15), .ZN(N7) );
  AOI22_X1 U5 ( .A1(port0[5]), .A2(n13), .B1(port1[5]), .B2(sel), .ZN(n15) );
  INV_X1 U6 ( .A(n20), .ZN(N2) );
  AOI22_X1 U7 ( .A1(port0[0]), .A2(n13), .B1(port1[0]), .B2(sel), .ZN(n20) );
  INV_X1 U8 ( .A(n19), .ZN(N3) );
  AOI22_X1 U9 ( .A1(port0[1]), .A2(n13), .B1(port1[1]), .B2(sel), .ZN(n19) );
  INV_X1 U10 ( .A(n18), .ZN(N4) );
  AOI22_X1 U11 ( .A1(port0[2]), .A2(n13), .B1(port1[2]), .B2(sel), .ZN(n18) );
  INV_X1 U12 ( .A(n17), .ZN(N5) );
  AOI22_X1 U13 ( .A1(port0[3]), .A2(n13), .B1(port1[3]), .B2(sel), .ZN(n17) );
  INV_X1 U14 ( .A(n12), .ZN(N9) );
  AOI22_X1 U15 ( .A1(port0[7]), .A2(n13), .B1(sel), .B2(port1[7]), .ZN(n12) );
  INV_X1 U16 ( .A(n21), .ZN(N11) );
  AOI22_X1 U17 ( .A1(port0[9]), .A2(n13), .B1(port1[9]), .B2(sel), .ZN(n21) );
  INV_X1 U18 ( .A(n14), .ZN(N8) );
  AOI22_X1 U19 ( .A1(port0[6]), .A2(n13), .B1(port1[6]), .B2(sel), .ZN(n14) );
  INV_X1 U20 ( .A(n22), .ZN(N10) );
  AOI22_X1 U21 ( .A1(port0[8]), .A2(n13), .B1(port1[8]), .B2(sel), .ZN(n22) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_79 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n5), .Z(n14) );
  BUF_X1 U4 ( .A(n4), .Z(n11) );
  BUF_X1 U5 ( .A(n4), .Z(n10) );
  BUF_X1 U6 ( .A(n6), .Z(n17) );
  BUF_X1 U7 ( .A(n4), .Z(n9) );
  BUF_X1 U8 ( .A(n6), .Z(n15) );
  BUF_X1 U9 ( .A(n6), .Z(n16) );
  BUF_X1 U10 ( .A(n5), .Z(n13) );
  BUF_X1 U11 ( .A(n5), .Z(n12) );
  BUF_X1 U12 ( .A(sel), .Z(n6) );
  BUF_X1 U13 ( .A(sel), .Z(n5) );
  BUF_X1 U14 ( .A(sel), .Z(n4) );
  INV_X1 U15 ( .A(n38), .ZN(N6) );
  INV_X1 U16 ( .A(n39), .ZN(N5) );
  INV_X1 U17 ( .A(n40), .ZN(N4) );
  INV_X1 U18 ( .A(n56), .ZN(N2) );
  INV_X1 U19 ( .A(n45), .ZN(N3) );
  INV_X1 U20 ( .A(n37), .ZN(N7) );
  INV_X1 U21 ( .A(n34), .ZN(N9) );
  INV_X1 U22 ( .A(n36), .ZN(N8) );
  INV_X1 U23 ( .A(n41), .ZN(N33) );
  INV_X1 U24 ( .A(n42), .ZN(N32) );
  INV_X1 U25 ( .A(n58), .ZN(N18) );
  INV_X1 U26 ( .A(n53), .ZN(N22) );
  INV_X1 U27 ( .A(n52), .ZN(N23) );
  INV_X1 U28 ( .A(n51), .ZN(N24) );
  INV_X1 U29 ( .A(n50), .ZN(N25) );
  INV_X1 U30 ( .A(n49), .ZN(N26) );
  INV_X1 U31 ( .A(n48), .ZN(N27) );
  INV_X1 U32 ( .A(n47), .ZN(N28) );
  INV_X1 U33 ( .A(n46), .ZN(N29) );
  INV_X1 U34 ( .A(n44), .ZN(N30) );
  INV_X1 U35 ( .A(n43), .ZN(N31) );
  INV_X1 U36 ( .A(n57), .ZN(N19) );
  INV_X1 U37 ( .A(n61), .ZN(N15) );
  INV_X1 U38 ( .A(n62), .ZN(N14) );
  INV_X1 U39 ( .A(n60), .ZN(N16) );
  INV_X1 U40 ( .A(n59), .ZN(N17) );
  INV_X1 U41 ( .A(n63), .ZN(N13) );
  INV_X1 U42 ( .A(n55), .ZN(N20) );
  INV_X1 U43 ( .A(n54), .ZN(N21) );
  INV_X1 U44 ( .A(n64), .ZN(N12) );
  INV_X1 U45 ( .A(n65), .ZN(N11) );
  INV_X1 U46 ( .A(n66), .ZN(N10) );
  AOI22_X1 U47 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n38) );
  AOI22_X1 U48 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n39) );
  AOI22_X1 U49 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(n10), .ZN(n40) );
  AOI22_X1 U50 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n56) );
  AOI22_X1 U51 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n45) );
  AOI22_X1 U52 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n37) );
  AOI22_X1 U53 ( .A1(port0[7]), .A2(n8), .B1(n16), .B2(port1[7]), .ZN(n34) );
  AOI22_X1 U54 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n36) );
  AOI22_X1 U55 ( .A1(port0[31]), .A2(n8), .B1(port1[31]), .B2(n10), .ZN(n41)
         );
  AOI22_X1 U56 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n42)
         );
  AOI22_X1 U57 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n57)
         );
  AOI22_X1 U58 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n64)
         );
  AOI22_X1 U59 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n61)
         );
  AOI22_X1 U60 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n62)
         );
  AOI22_X1 U61 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n60)
         );
  AOI22_X1 U62 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n65) );
  AOI22_X1 U63 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n66) );
  AOI22_X1 U64 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n59)
         );
  AOI22_X1 U65 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n63)
         );
  AOI22_X1 U66 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n58)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n55)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n54)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n53)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n52)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n51)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n49)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n48)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n47)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n46)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n44)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n43)
         );
endmodule


module Enable_Interface_NBIT_DATA5_0 ( EI_datain, EI_enable, EI_dataout );
  input [4:0] EI_datain;
  output [4:0] EI_dataout;
  input EI_enable;


  AND2_X1 U1 ( .A1(EI_datain[3]), .A2(EI_enable), .ZN(EI_dataout[3]) );
  AND2_X1 U2 ( .A1(EI_datain[0]), .A2(EI_enable), .ZN(EI_dataout[0]) );
  AND2_X1 U3 ( .A1(EI_enable), .A2(EI_datain[4]), .ZN(EI_dataout[4]) );
  AND2_X1 U4 ( .A1(EI_datain[1]), .A2(EI_enable), .ZN(EI_dataout[1]) );
  AND2_X1 U5 ( .A1(EI_datain[2]), .A2(EI_enable), .ZN(EI_dataout[2]) );
endmodule


module Decoder_DEC_NBIT5 ( DEC_address, DEC_enable, DEC_output );
  input [4:0] DEC_address;
  output [31:0] DEC_output;
  input DEC_enable;
  wire   n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20,
         n21, n22;

  NAND3_X1 U39 ( .A1(DEC_enable), .A2(DEC_address[3]), .A3(DEC_address[4]), 
        .ZN(n15) );
  NAND3_X1 U40 ( .A1(n18), .A2(n19), .A3(DEC_address[0]), .ZN(n6) );
  NAND3_X1 U41 ( .A1(DEC_enable), .A2(n20), .A3(DEC_address[4]), .ZN(n17) );
  NAND3_X1 U42 ( .A1(DEC_address[1]), .A2(DEC_address[0]), .A3(DEC_address[2]), 
        .ZN(n9) );
  NAND3_X1 U43 ( .A1(DEC_address[1]), .A2(n21), .A3(DEC_address[2]), .ZN(n11)
         );
  NAND3_X1 U44 ( .A1(DEC_address[0]), .A2(n18), .A3(DEC_address[2]), .ZN(n12)
         );
  NAND3_X1 U45 ( .A1(n21), .A2(n18), .A3(DEC_address[2]), .ZN(n13) );
  NAND3_X1 U46 ( .A1(DEC_address[0]), .A2(n19), .A3(DEC_address[1]), .ZN(n14)
         );
  NAND3_X1 U47 ( .A1(n21), .A2(n19), .A3(DEC_address[1]), .ZN(n16) );
  NAND3_X1 U48 ( .A1(DEC_address[3]), .A2(n22), .A3(DEC_enable), .ZN(n7) );
  NAND3_X1 U49 ( .A1(n20), .A2(n22), .A3(DEC_enable), .ZN(n10) );
  NAND3_X1 U50 ( .A1(n18), .A2(n19), .A3(n21), .ZN(n8) );
  NOR2_X1 U2 ( .A1(n8), .A2(n10), .ZN(DEC_output[0]) );
  NOR2_X1 U3 ( .A1(n10), .A2(n16), .ZN(DEC_output[2]) );
  NOR2_X1 U4 ( .A1(n10), .A2(n14), .ZN(DEC_output[3]) );
  NOR2_X1 U5 ( .A1(n10), .A2(n13), .ZN(DEC_output[4]) );
  NOR2_X1 U6 ( .A1(n10), .A2(n12), .ZN(DEC_output[5]) );
  NOR2_X1 U7 ( .A1(n10), .A2(n11), .ZN(DEC_output[6]) );
  NOR2_X1 U8 ( .A1(n9), .A2(n10), .ZN(DEC_output[7]) );
  NOR2_X1 U9 ( .A1(n6), .A2(n7), .ZN(DEC_output[9]) );
  NOR2_X1 U10 ( .A1(n7), .A2(n16), .ZN(DEC_output[10]) );
  NOR2_X1 U11 ( .A1(n7), .A2(n14), .ZN(DEC_output[11]) );
  NOR2_X1 U12 ( .A1(n7), .A2(n13), .ZN(DEC_output[12]) );
  NOR2_X1 U13 ( .A1(n7), .A2(n12), .ZN(DEC_output[13]) );
  NOR2_X1 U14 ( .A1(n7), .A2(n11), .ZN(DEC_output[14]) );
  NOR2_X1 U15 ( .A1(n7), .A2(n9), .ZN(DEC_output[15]) );
  NOR2_X1 U16 ( .A1(n8), .A2(n17), .ZN(DEC_output[16]) );
  NOR2_X1 U17 ( .A1(n6), .A2(n17), .ZN(DEC_output[17]) );
  NOR2_X1 U18 ( .A1(n14), .A2(n17), .ZN(DEC_output[19]) );
  NOR2_X1 U19 ( .A1(n13), .A2(n17), .ZN(DEC_output[20]) );
  NOR2_X1 U20 ( .A1(n12), .A2(n17), .ZN(DEC_output[21]) );
  NOR2_X1 U21 ( .A1(n11), .A2(n17), .ZN(DEC_output[22]) );
  NOR2_X1 U22 ( .A1(n9), .A2(n17), .ZN(DEC_output[23]) );
  NOR2_X1 U23 ( .A1(n8), .A2(n15), .ZN(DEC_output[24]) );
  NOR2_X1 U24 ( .A1(n6), .A2(n15), .ZN(DEC_output[25]) );
  NOR2_X1 U25 ( .A1(n15), .A2(n16), .ZN(DEC_output[26]) );
  NOR2_X1 U26 ( .A1(n13), .A2(n15), .ZN(DEC_output[28]) );
  NOR2_X1 U27 ( .A1(n12), .A2(n15), .ZN(DEC_output[29]) );
  NOR2_X1 U28 ( .A1(n11), .A2(n15), .ZN(DEC_output[30]) );
  NOR2_X1 U29 ( .A1(n9), .A2(n15), .ZN(DEC_output[31]) );
  NOR2_X1 U30 ( .A1(n6), .A2(n10), .ZN(DEC_output[1]) );
  NOR2_X1 U31 ( .A1(n7), .A2(n8), .ZN(DEC_output[8]) );
  NOR2_X1 U32 ( .A1(n16), .A2(n17), .ZN(DEC_output[18]) );
  NOR2_X1 U33 ( .A1(n14), .A2(n15), .ZN(DEC_output[27]) );
  INV_X1 U34 ( .A(DEC_address[2]), .ZN(n19) );
  INV_X1 U35 ( .A(DEC_address[0]), .ZN(n21) );
  INV_X1 U36 ( .A(DEC_address[1]), .ZN(n18) );
  INV_X1 U37 ( .A(DEC_address[4]), .ZN(n22) );
  INV_X1 U38 ( .A(DEC_address[3]), .ZN(n20) );
endmodule


module Sum_Network_N32_0 ( G, P, S );
  input [31:0] G;
  input [31:0] P;
  output [31:0] S;


  XOR2_X1 U1 ( .A(P[9]), .B(G[9]), .Z(S[9]) );
  XOR2_X1 U2 ( .A(P[8]), .B(G[8]), .Z(S[8]) );
  XOR2_X1 U3 ( .A(P[7]), .B(G[7]), .Z(S[7]) );
  XOR2_X1 U4 ( .A(P[6]), .B(G[6]), .Z(S[6]) );
  XOR2_X1 U5 ( .A(P[5]), .B(G[5]), .Z(S[5]) );
  XOR2_X1 U6 ( .A(P[4]), .B(G[4]), .Z(S[4]) );
  XOR2_X1 U7 ( .A(P[3]), .B(G[3]), .Z(S[3]) );
  XOR2_X1 U8 ( .A(P[31]), .B(G[31]), .Z(S[31]) );
  XOR2_X1 U9 ( .A(P[30]), .B(G[30]), .Z(S[30]) );
  XOR2_X1 U10 ( .A(P[2]), .B(G[2]), .Z(S[2]) );
  XOR2_X1 U11 ( .A(P[29]), .B(G[29]), .Z(S[29]) );
  XOR2_X1 U12 ( .A(P[28]), .B(G[28]), .Z(S[28]) );
  XOR2_X1 U13 ( .A(P[27]), .B(G[27]), .Z(S[27]) );
  XOR2_X1 U14 ( .A(P[26]), .B(G[26]), .Z(S[26]) );
  XOR2_X1 U15 ( .A(P[25]), .B(G[25]), .Z(S[25]) );
  XOR2_X1 U16 ( .A(P[24]), .B(G[24]), .Z(S[24]) );
  XOR2_X1 U17 ( .A(P[23]), .B(G[23]), .Z(S[23]) );
  XOR2_X1 U18 ( .A(P[22]), .B(G[22]), .Z(S[22]) );
  XOR2_X1 U19 ( .A(P[21]), .B(G[21]), .Z(S[21]) );
  XOR2_X1 U20 ( .A(P[20]), .B(G[20]), .Z(S[20]) );
  XOR2_X1 U21 ( .A(P[1]), .B(G[1]), .Z(S[1]) );
  XOR2_X1 U22 ( .A(P[19]), .B(G[19]), .Z(S[19]) );
  XOR2_X1 U23 ( .A(P[18]), .B(G[18]), .Z(S[18]) );
  XOR2_X1 U24 ( .A(P[17]), .B(G[17]), .Z(S[17]) );
  XOR2_X1 U25 ( .A(P[16]), .B(G[16]), .Z(S[16]) );
  XOR2_X1 U26 ( .A(P[15]), .B(G[15]), .Z(S[15]) );
  XOR2_X1 U27 ( .A(P[14]), .B(G[14]), .Z(S[14]) );
  XOR2_X1 U28 ( .A(P[13]), .B(G[13]), .Z(S[13]) );
  XOR2_X1 U29 ( .A(P[12]), .B(G[12]), .Z(S[12]) );
  XOR2_X1 U30 ( .A(P[11]), .B(G[11]), .Z(S[11]) );
  XOR2_X1 U31 ( .A(P[10]), .B(G[10]), .Z(S[10]) );
  XOR2_X1 U32 ( .A(P[0]), .B(G[0]), .Z(S[0]) );
endmodule


module Carry_Network_N32_0 ( G, P, Cin, Cout, Gout, Pout );
  input [31:0] G;
  input [31:0] P;
  output [31:0] Gout;
  output [31:0] Pout;
  input Cin;
  output Cout;
  wire   Cin, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64;
  assign Gout[0] = Cin;
  assign Pout[31] = P[31];
  assign Pout[30] = P[30];
  assign Pout[29] = P[29];
  assign Pout[28] = P[28];
  assign Pout[27] = P[27];
  assign Pout[26] = P[26];
  assign Pout[25] = P[25];
  assign Pout[24] = P[24];
  assign Pout[23] = P[23];
  assign Pout[22] = P[22];
  assign Pout[21] = P[21];
  assign Pout[20] = P[20];
  assign Pout[19] = P[19];
  assign Pout[18] = P[18];
  assign Pout[17] = P[17];
  assign Pout[16] = P[16];
  assign Pout[15] = P[15];
  assign Pout[14] = P[14];
  assign Pout[13] = P[13];
  assign Pout[12] = P[12];
  assign Pout[11] = P[11];
  assign Pout[10] = P[10];
  assign Pout[9] = P[9];
  assign Pout[8] = P[8];
  assign Pout[7] = P[7];
  assign Pout[6] = P[6];
  assign Pout[5] = P[5];
  assign Pout[4] = P[4];
  assign Pout[3] = P[3];
  assign Pout[2] = P[2];
  assign Pout[1] = P[1];
  assign Pout[0] = P[0];

  INV_X1 U1 ( .A(n33), .ZN(Cout) );
  INV_X1 U2 ( .A(n63), .ZN(Gout[2]) );
  AOI21_X1 U3 ( .B1(P[1]), .B2(Gout[1]), .A(G[1]), .ZN(n63) );
  INV_X1 U4 ( .A(n62), .ZN(Gout[3]) );
  AOI21_X1 U5 ( .B1(P[2]), .B2(Gout[2]), .A(G[2]), .ZN(n62) );
  INV_X1 U6 ( .A(n61), .ZN(Gout[4]) );
  AOI21_X1 U7 ( .B1(P[3]), .B2(Gout[3]), .A(G[3]), .ZN(n61) );
  INV_X1 U8 ( .A(n60), .ZN(Gout[5]) );
  AOI21_X1 U9 ( .B1(P[4]), .B2(Gout[4]), .A(G[4]), .ZN(n60) );
  INV_X1 U10 ( .A(n59), .ZN(Gout[6]) );
  AOI21_X1 U11 ( .B1(P[5]), .B2(Gout[5]), .A(G[5]), .ZN(n59) );
  INV_X1 U12 ( .A(n58), .ZN(Gout[7]) );
  AOI21_X1 U13 ( .B1(P[6]), .B2(Gout[6]), .A(G[6]), .ZN(n58) );
  INV_X1 U14 ( .A(n57), .ZN(Gout[8]) );
  AOI21_X1 U15 ( .B1(P[7]), .B2(Gout[7]), .A(G[7]), .ZN(n57) );
  INV_X1 U16 ( .A(n56), .ZN(Gout[9]) );
  AOI21_X1 U17 ( .B1(P[8]), .B2(Gout[8]), .A(G[8]), .ZN(n56) );
  INV_X1 U18 ( .A(n55), .ZN(Gout[10]) );
  AOI21_X1 U19 ( .B1(P[9]), .B2(Gout[9]), .A(G[9]), .ZN(n55) );
  INV_X1 U20 ( .A(n54), .ZN(Gout[11]) );
  AOI21_X1 U21 ( .B1(P[10]), .B2(Gout[10]), .A(G[10]), .ZN(n54) );
  INV_X1 U22 ( .A(n53), .ZN(Gout[12]) );
  AOI21_X1 U23 ( .B1(P[11]), .B2(Gout[11]), .A(G[11]), .ZN(n53) );
  INV_X1 U24 ( .A(n52), .ZN(Gout[13]) );
  AOI21_X1 U25 ( .B1(P[12]), .B2(Gout[12]), .A(G[12]), .ZN(n52) );
  INV_X1 U26 ( .A(n51), .ZN(Gout[14]) );
  AOI21_X1 U27 ( .B1(P[13]), .B2(Gout[13]), .A(G[13]), .ZN(n51) );
  INV_X1 U28 ( .A(n50), .ZN(Gout[15]) );
  AOI21_X1 U29 ( .B1(P[14]), .B2(Gout[14]), .A(G[14]), .ZN(n50) );
  INV_X1 U30 ( .A(n49), .ZN(Gout[16]) );
  AOI21_X1 U31 ( .B1(P[15]), .B2(Gout[15]), .A(G[15]), .ZN(n49) );
  INV_X1 U32 ( .A(n48), .ZN(Gout[17]) );
  AOI21_X1 U33 ( .B1(P[16]), .B2(Gout[16]), .A(G[16]), .ZN(n48) );
  INV_X1 U34 ( .A(n47), .ZN(Gout[18]) );
  AOI21_X1 U35 ( .B1(P[17]), .B2(Gout[17]), .A(G[17]), .ZN(n47) );
  INV_X1 U36 ( .A(n46), .ZN(Gout[19]) );
  AOI21_X1 U37 ( .B1(P[18]), .B2(Gout[18]), .A(G[18]), .ZN(n46) );
  INV_X1 U38 ( .A(n45), .ZN(Gout[20]) );
  AOI21_X1 U39 ( .B1(P[19]), .B2(Gout[19]), .A(G[19]), .ZN(n45) );
  INV_X1 U40 ( .A(n44), .ZN(Gout[21]) );
  AOI21_X1 U41 ( .B1(P[20]), .B2(Gout[20]), .A(G[20]), .ZN(n44) );
  INV_X1 U42 ( .A(n43), .ZN(Gout[22]) );
  AOI21_X1 U43 ( .B1(P[21]), .B2(Gout[21]), .A(G[21]), .ZN(n43) );
  INV_X1 U44 ( .A(n42), .ZN(Gout[23]) );
  AOI21_X1 U45 ( .B1(P[22]), .B2(Gout[22]), .A(G[22]), .ZN(n42) );
  INV_X1 U46 ( .A(n41), .ZN(Gout[24]) );
  AOI21_X1 U47 ( .B1(P[23]), .B2(Gout[23]), .A(G[23]), .ZN(n41) );
  INV_X1 U48 ( .A(n40), .ZN(Gout[25]) );
  AOI21_X1 U49 ( .B1(P[24]), .B2(Gout[24]), .A(G[24]), .ZN(n40) );
  INV_X1 U50 ( .A(n39), .ZN(Gout[26]) );
  AOI21_X1 U51 ( .B1(P[25]), .B2(Gout[25]), .A(G[25]), .ZN(n39) );
  INV_X1 U52 ( .A(n38), .ZN(Gout[27]) );
  AOI21_X1 U53 ( .B1(P[26]), .B2(Gout[26]), .A(G[26]), .ZN(n38) );
  INV_X1 U54 ( .A(n37), .ZN(Gout[28]) );
  AOI21_X1 U55 ( .B1(P[27]), .B2(Gout[27]), .A(G[27]), .ZN(n37) );
  INV_X1 U56 ( .A(n36), .ZN(Gout[29]) );
  AOI21_X1 U57 ( .B1(P[28]), .B2(Gout[28]), .A(G[28]), .ZN(n36) );
  INV_X1 U58 ( .A(n35), .ZN(Gout[30]) );
  AOI21_X1 U59 ( .B1(P[29]), .B2(Gout[29]), .A(G[29]), .ZN(n35) );
  INV_X1 U60 ( .A(n34), .ZN(Gout[31]) );
  AOI21_X1 U61 ( .B1(P[30]), .B2(Gout[30]), .A(G[30]), .ZN(n34) );
  INV_X1 U62 ( .A(n64), .ZN(Gout[1]) );
  AOI21_X1 U63 ( .B1(P[0]), .B2(Cin), .A(G[0]), .ZN(n64) );
  AOI21_X1 U64 ( .B1(P[31]), .B2(Gout[31]), .A(G[31]), .ZN(n33) );
endmodule


module PG_network_N32_0 ( A, B, c_in, G, P );
  input [31:0] A;
  input [31:0] B;
  output [31:0] G;
  output [31:0] P;
  input c_in;
  wire   tmp1, tmp2;
  assign P[0] = 1'b0;

  XOR2_X1 U3 ( .A(B[0]), .B(A[0]), .Z(tmp2) );
  GeneralGenerate_0 G_cell_0_0 ( .G_ik(tmp1), .P_ik(tmp2), .G_km1_j(c_in), 
        .G_ij(G[0]) );
  PG_cell_0 PG_cell_i_1 ( .A(A[1]), .B(B[1]), .p(P[1]), .g(G[1]) );
  PG_cell_92 PG_cell_i_2 ( .A(A[2]), .B(B[2]), .p(P[2]), .g(G[2]) );
  PG_cell_91 PG_cell_i_3 ( .A(A[3]), .B(B[3]), .p(P[3]), .g(G[3]) );
  PG_cell_90 PG_cell_i_4 ( .A(A[4]), .B(B[4]), .p(P[4]), .g(G[4]) );
  PG_cell_89 PG_cell_i_5 ( .A(A[5]), .B(B[5]), .p(P[5]), .g(G[5]) );
  PG_cell_88 PG_cell_i_6 ( .A(A[6]), .B(B[6]), .p(P[6]), .g(G[6]) );
  PG_cell_87 PG_cell_i_7 ( .A(A[7]), .B(B[7]), .p(P[7]), .g(G[7]) );
  PG_cell_86 PG_cell_i_8 ( .A(A[8]), .B(B[8]), .p(P[8]), .g(G[8]) );
  PG_cell_85 PG_cell_i_9 ( .A(A[9]), .B(B[9]), .p(P[9]), .g(G[9]) );
  PG_cell_84 PG_cell_i_10 ( .A(A[10]), .B(B[10]), .p(P[10]), .g(G[10]) );
  PG_cell_83 PG_cell_i_11 ( .A(A[11]), .B(B[11]), .p(P[11]), .g(G[11]) );
  PG_cell_82 PG_cell_i_12 ( .A(A[12]), .B(B[12]), .p(P[12]), .g(G[12]) );
  PG_cell_81 PG_cell_i_13 ( .A(A[13]), .B(B[13]), .p(P[13]), .g(G[13]) );
  PG_cell_80 PG_cell_i_14 ( .A(A[14]), .B(B[14]), .p(P[14]), .g(G[14]) );
  PG_cell_79 PG_cell_i_15 ( .A(A[15]), .B(B[15]), .p(P[15]), .g(G[15]) );
  PG_cell_78 PG_cell_i_16 ( .A(A[16]), .B(B[16]), .p(P[16]), .g(G[16]) );
  PG_cell_77 PG_cell_i_17 ( .A(A[17]), .B(B[17]), .p(P[17]), .g(G[17]) );
  PG_cell_76 PG_cell_i_18 ( .A(A[18]), .B(B[18]), .p(P[18]), .g(G[18]) );
  PG_cell_75 PG_cell_i_19 ( .A(A[19]), .B(B[19]), .p(P[19]), .g(G[19]) );
  PG_cell_74 PG_cell_i_20 ( .A(A[20]), .B(B[20]), .p(P[20]), .g(G[20]) );
  PG_cell_73 PG_cell_i_21 ( .A(A[21]), .B(B[21]), .p(P[21]), .g(G[21]) );
  PG_cell_72 PG_cell_i_22 ( .A(A[22]), .B(B[22]), .p(P[22]), .g(G[22]) );
  PG_cell_71 PG_cell_i_23 ( .A(A[23]), .B(B[23]), .p(P[23]), .g(G[23]) );
  PG_cell_70 PG_cell_i_24 ( .A(A[24]), .B(B[24]), .p(P[24]), .g(G[24]) );
  PG_cell_69 PG_cell_i_25 ( .A(A[25]), .B(B[25]), .p(P[25]), .g(G[25]) );
  PG_cell_68 PG_cell_i_26 ( .A(A[26]), .B(B[26]), .p(P[26]), .g(G[26]) );
  PG_cell_67 PG_cell_i_27 ( .A(A[27]), .B(B[27]), .p(P[27]), .g(G[27]) );
  PG_cell_66 PG_cell_i_28 ( .A(A[28]), .B(B[28]), .p(P[28]), .g(G[28]) );
  PG_cell_65 PG_cell_i_29 ( .A(A[29]), .B(B[29]), .p(P[29]), .g(G[29]) );
  PG_cell_64 PG_cell_i_30 ( .A(A[30]), .B(B[30]), .p(P[30]), .g(G[30]) );
  PG_cell_63 PG_cell_i_31 ( .A(A[31]), .B(B[31]), .p(P[31]), .g(G[31]) );
  AND2_X1 U2 ( .A1(B[0]), .A2(A[0]), .ZN(tmp1) );
endmodule


module UD_COUNTER_BTB_UDC_NBIT3_0 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT
 );
  output [2:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   n3, n5, n6;
  wire   [1:0] s_nq;
  wire   [2:1] s_toggle;

  NAND3_X1 U5 ( .A1(UDC_OUT[0]), .A2(UDC_EN), .A3(UDC_UP), .ZN(n5) );
  NAND3_X1 U6 ( .A1(UDC_EN), .A2(n6), .A3(s_nq[0]), .ZN(n3) );
  t_ff_rst0_64 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(s_nq[0]) );
  t_ff_rst0_63 FF_i_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[1]), .TFF_q(UDC_OUT[1]), .TFF_nq(s_nq[1]) );
  t_ff_rst1_32 FF_N_2 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        s_toggle[2]), .TFF_q(UDC_OUT[2]) );
  OAI22_X1 U1 ( .A1(n3), .A2(UDC_OUT[1]), .B1(s_nq[1]), .B2(n5), .ZN(
        s_toggle[2]) );
  INV_X1 U2 ( .A(UDC_UP), .ZN(n6) );
  NAND2_X1 U3 ( .A1(n3), .A2(n5), .ZN(s_toggle[1]) );
endmodule


module Mux_Bit_NBIT_Sel2_0 ( inputs, sel, \output  );
  input [3:0] inputs;
  input [1:0] sel;
  output \output ;
  wire   n3, n5, n4, n6;

  OAI22_X1 U1 ( .A1(n3), .A2(n6), .B1(sel[1]), .B2(n5), .ZN(\output ) );
  AOI22_X1 U2 ( .A1(inputs[2]), .A2(n4), .B1(inputs[3]), .B2(sel[0]), .ZN(n3)
         );
  AOI22_X1 U3 ( .A1(inputs[0]), .A2(n4), .B1(sel[0]), .B2(inputs[1]), .ZN(n5)
         );
  INV_X1 U4 ( .A(sel[0]), .ZN(n4) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n6) );
endmodule


module D_FF_0 ( D, clk, Q, Not_Q );
  input D, clk;
  output Q, Not_Q;
  wire   N0;

  DFF_X1 Q_reg ( .D(D), .CK(clk), .Q(Q) );
  DFF_X1 Not_Q_reg ( .D(N0), .CK(clk), .Q(Not_Q) );
  INV_X1 U3 ( .A(D), .ZN(N0) );
endmodule


module ComparatorWithEnable_0 ( a, b, enable, y );
  input a, b, enable;
  output y;
  wire   n1;

  AND2_X1 U1 ( .A1(n1), .A2(enable), .ZN(y) );
  XNOR2_X1 U2 ( .A(b), .B(a), .ZN(n1) );
endmodule


module NORGate_NX1_N2 ( A, B, Y );
  input [1:0] A;
  input [1:0] B;
  output Y;


  NOR4_X1 U1 ( .A1(B[1]), .A2(B[0]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module ANDGate_NX1_N2 ( A, B, Y );
  input [1:0] A;
  input [1:0] B;
  output Y;


  AND4_X1 U1 ( .A1(B[1]), .A2(B[0]), .A3(A[1]), .A4(A[0]), .ZN(Y) );
endmodule


module CU_SatCounter_0 ( CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, 
        CU_loadDefault, CU_TcMax, CU_TcMin, UDC_clk, UDC_Ud, UDC_enable, 
        UDC_reset );
  input CU_clk, CU_reset, CU_enable, CU_Ud, CU_update, CU_loadDefault,
         CU_TcMax, CU_TcMin;
  output UDC_clk, UDC_Ud, UDC_enable, UDC_reset;
  wire   CU_clk, n5, n6, n7, n8, n9, n10;
  assign UDC_clk = CU_clk;

  NOR3_X1 U3 ( .A1(CU_TcMax), .A2(n7), .A3(n8), .ZN(UDC_Ud) );
  INV_X1 U4 ( .A(CU_Ud), .ZN(n8) );
  NAND4_X1 U5 ( .A1(CU_update), .A2(CU_enable), .A3(n9), .A4(n10), .ZN(n7) );
  INV_X1 U6 ( .A(CU_loadDefault), .ZN(n9) );
  OR2_X1 U7 ( .A1(n6), .A2(UDC_Ud), .ZN(UDC_enable) );
  NOR3_X1 U8 ( .A1(n7), .A2(CU_Ud), .A3(CU_TcMin), .ZN(n6) );
  INV_X1 U9 ( .A(n5), .ZN(UDC_reset) );
  AOI21_X1 U10 ( .B1(CU_enable), .B2(CU_loadDefault), .A(CU_reset), .ZN(n5) );
  INV_X1 U11 ( .A(CU_reset), .ZN(n10) );
endmodule


module UD_COUNTER_UDC_NBIT2 ( UDC_EN, UDC_UP, UDC_CLK, UDC_RST, UDC_OUT );
  output [1:0] UDC_OUT;
  input UDC_EN, UDC_UP, UDC_CLK, UDC_RST;
  wire   \s_nq[0] , \s_toggle[1] , n1;

  XOR2_X1 U2 ( .A(\s_nq[0] ), .B(UDC_UP), .Z(n1) );
  t_ff_rst1_0 FF_0_0 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(UDC_EN), 
        .TFF_q(UDC_OUT[0]), .TFF_nq(\s_nq[0] ) );
  t_ff_rst0_0 FF_N_1 ( .TFF_clk(UDC_CLK), .TFF_rst(UDC_RST), .TFF_t(
        \s_toggle[1] ), .TFF_q(UDC_OUT[1]) );
  AND2_X1 U1 ( .A1(UDC_EN), .A2(n1), .ZN(\s_toggle[1] ) );
endmodule


module Sign_Reducer_NBIT_data32 ( SR_data_in, SR_reduce, SR_BYTE_half, 
        SR_SGN_usg, SR_data_out );
  input [31:0] SR_data_in;
  output [31:0] SR_data_out;
  input SR_reduce, SR_BYTE_half, SR_SGN_usg;
  wire   s_msb, \s_tmp[9] , n1, n2, n3, n4, n5, n6, n7, n8, n9;
  wire   [31:0] s_tmp2;

  Mux_1Bit_2X1_3 MUX_msb ( .port0(SR_data_in[15]), .port1(SR_data_in[7]), 
        .sel(SR_BYTE_half), .portY(s_msb) );
  Mux_NBit_2x1_NBIT_IN32_9 MUX_B_H ( .port0({n3, n5, n5, n2, n2, n7, n3, n3, 
        n2, n3, n1, n3, n2, n7, n3, n3, n6, SR_data_in[14:8], n8, 
        SR_data_in[6:0]}), .port1({n2, \s_tmp[9] , \s_tmp[9] , n7, n5, n3, n2, 
        n5, n7, n7, n7, n7, n2, n3, n1, n7, n3, n7, n3, n3, n7, n7, n3, n7, n8, 
        SR_data_in[6:0]}), .sel(SR_BYTE_half), .portY(s_tmp2) );
  Mux_NBit_2x1_NBIT_IN32_8 MUX_OUT ( .port0({SR_data_in[31:16], n6, 
        SR_data_in[14:8], n9, SR_data_in[6:2], n4, SR_data_in[0]}), .port1(
        s_tmp2), .sel(SR_reduce), .portY(SR_data_out) );
  CLKBUF_X1 U1 ( .A(\s_tmp[9] ), .Z(n1) );
  AND2_X1 U2 ( .A1(s_msb), .A2(SR_SGN_usg), .ZN(\s_tmp[9] ) );
  AND2_X1 U3 ( .A1(s_msb), .A2(SR_SGN_usg), .ZN(n2) );
  AND2_X2 U4 ( .A1(s_msb), .A2(SR_SGN_usg), .ZN(n3) );
  AND2_X1 U5 ( .A1(s_msb), .A2(SR_SGN_usg), .ZN(n5) );
  CLKBUF_X1 U6 ( .A(SR_data_in[1]), .Z(n4) );
  AND2_X2 U7 ( .A1(s_msb), .A2(SR_SGN_usg), .ZN(n7) );
  CLKBUF_X1 U8 ( .A(SR_data_in[15]), .Z(n6) );
  CLKBUF_X1 U9 ( .A(SR_data_in[7]), .Z(n8) );
  CLKBUF_X1 U10 ( .A(n8), .Z(n9) );
endmodule


module Data_Reducer_NBIT_DATA32 ( DR_data_in, DR_reduce, DR_BYTE_half, 
        DR_data_out );
  input [31:0] DR_data_in;
  output [31:0] DR_data_out;
  input DR_reduce, DR_BYTE_half;

  wire   [31:0] s_tmp;

  Mux_NBit_2x1_NBIT_IN32_11 MUX_B_H ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        DR_data_in[15:0]}), .port1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, DR_data_in[7:0]}), .sel(DR_BYTE_half), 
        .portY(s_tmp) );
  Mux_NBit_2x1_NBIT_IN32_10 MUX_OUT ( .port0(DR_data_in), .port1(s_tmp), .sel(
        DR_reduce), .portY(DR_data_out) );
endmodule


module Multiplier_NBIT_DATA32 ( MUL_OpA, MUL_OpB, MUL_SGN_usgn, MUL_product );
  input [31:0] MUL_OpA;
  input [31:0] MUL_OpB;
  output [63:0] MUL_product;
  input MUL_SGN_usgn;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, N34, N35, N36, N37, N38, N39, N40, N41, N42, N43, N44,
         N45, N46, N47, N48, N49, N50, N51, N52, N53, N54, N55, N56, N57, N58,
         N59, N60, N61, N62, N63, N64, N65, N66, N67, N68, N69, N70, N71, N72,
         N73, N74, N75, N76, N77, N78, N79, N80, N81, N82, N83, N84, N85, N86,
         N87, N88, N89, N90, N91, N92, N93, N94, N95, N96, N97, N98, N99, N100,
         N101, N102, N103, N104, N105, N106, N107, N108, N109, N110, N111,
         N112, N113, N114, N115, N116, N117, N118, N119, N120, N121, N122,
         N123, N124, N125, N126, N127, N128, N129, N130, N131, N132, N133,
         N134, N135, N136, N137, N138, N139, N140, N141, N142, N143, N144,
         N145, N146, N147, N148, N149, N150, N151, N152, N153, N154, N155,
         N156, N157, N158, N159, N160, N161, N162, N163, N164, N165, N166,
         N167, N168, N169, N170, N171, N172, N173, N174, N175, N176, N177,
         N178, N179, N180, N181, N182, N183, N184, N185, N186, N187, N188,
         N189, N190, N191, N192, N193, n72, n73, n74, n75, n76, n77, n78, n79,
         n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93,
         n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104, n105,
         n106, n107, n108, n109, n110, n111, n112, n113, n114, n115, n116,
         n117, n118, n119, n120, n121, n122, n123, n124, n125, n126, n127,
         n128, n129, n130, n131, n132, n133, n134, net132725, net132723,
         net132721, net132719, net132717, net132715, net132713, net132711,
         net132709, net132707, net132705, net132703, net132701, net132699,
         net132697, net132695, net132689, net132687, net132681, net132735,
         net132733, net132731, net132729, n3, n4, n5, n6, n7, n8, n9;
  assign MUL_product[0] = N130;
  assign MUL_product[1] = N131;
  assign MUL_product[2] = N132;
  assign MUL_product[3] = N133;
  assign MUL_product[4] = N134;
  assign MUL_product[5] = N135;
  assign MUL_product[6] = N136;
  assign MUL_product[7] = N137;
  assign MUL_product[8] = N138;
  assign MUL_product[9] = N139;
  assign MUL_product[10] = N140;
  assign MUL_product[11] = N141;
  assign MUL_product[12] = N142;
  assign MUL_product[13] = N143;
  assign MUL_product[14] = N144;
  assign MUL_product[15] = N145;
  assign MUL_product[16] = N146;
  assign MUL_product[17] = N147;
  assign MUL_product[18] = N148;
  assign MUL_product[19] = N149;
  assign MUL_product[20] = N150;
  assign MUL_product[21] = N151;
  assign MUL_product[22] = N152;
  assign MUL_product[23] = N153;
  assign MUL_product[24] = N154;
  assign MUL_product[25] = N155;
  assign MUL_product[26] = N156;
  assign MUL_product[27] = N157;
  assign MUL_product[28] = N158;
  assign MUL_product[29] = N159;
  assign MUL_product[30] = N160;
  assign MUL_product[31] = N161;
  assign MUL_product[32] = N162;
  assign MUL_product[33] = N163;
  assign MUL_product[34] = N164;
  assign MUL_product[35] = N165;
  assign MUL_product[36] = N166;
  assign MUL_product[37] = N167;
  assign MUL_product[38] = N168;
  assign MUL_product[39] = N169;
  assign MUL_product[40] = N170;
  assign MUL_product[41] = N171;
  assign MUL_product[42] = N172;
  assign MUL_product[43] = N173;
  assign MUL_product[44] = N174;
  assign MUL_product[45] = N175;
  assign MUL_product[46] = N176;
  assign MUL_product[47] = N177;
  assign MUL_product[48] = N178;
  assign MUL_product[49] = N179;
  assign MUL_product[50] = N180;
  assign MUL_product[51] = N181;
  assign MUL_product[52] = N182;
  assign MUL_product[53] = N183;
  assign MUL_product[54] = N184;
  assign MUL_product[55] = N185;
  assign MUL_product[56] = N186;
  assign MUL_product[57] = N187;
  assign MUL_product[58] = N188;
  assign MUL_product[59] = N189;
  assign MUL_product[60] = N190;
  assign MUL_product[61] = N191;
  assign MUL_product[62] = N192;
  assign MUL_product[63] = N193;

  Multiplier_NBIT_DATA32_DW02_mult_0 mult_65 ( .A(MUL_OpA), .B(MUL_OpB), .TC(
        1'b0), .PRODUCT({N129, N128, N127, N126, N125, N124, N123, N122, N121, 
        N120, N119, N118, N117, N116, N115, N114, N113, N112, N111, N110, N109, 
        N108, N107, N106, N105, N104, N103, N102, N101, N100, N99, N98, N97, 
        N96, N95, N94, N93, N92, N91, N90, N89, N88, N87, N86, N85, N84, N83, 
        N82, N81, N80, N79, N78, N77, N76, N75, N74, N73, N72, N71, N70, N69, 
        N68, N67, N66}) );
  Multiplier_NBIT_DATA32_DW02_mult_1 mult_61 ( .A(MUL_OpA), .B(MUL_OpB), .TC(
        1'b1), .PRODUCT({N65, N64, N63, N62, N61, N60, N59, N58, N57, N56, N55, 
        N54, N53, N52, N51, N50, N49, N48, N47, N46, N45, N44, N43, N42, N41, 
        N40, N39, N38, N37, N36, N35, N34, N33, N32, N31, N30, N29, N28, N27, 
        N26, N25, N24, N23, N22, N21, N20, N19, N18, N17, N16, N15, N14, N13, 
        N12, N11, N10, N9, N8, N7, N6, N5, N4, N3, N2}) );
  NAND2_X1 U1 ( .A1(N129), .A2(net132687), .ZN(n3) );
  NAND2_X1 U2 ( .A1(N65), .A2(net132723), .ZN(n4) );
  NAND2_X1 U5 ( .A1(n3), .A2(n4), .ZN(N193) );
  BUF_X1 U6 ( .A(n6), .Z(n5) );
  AOI22_X1 U7 ( .A1(N128), .A2(net132689), .B1(N64), .B2(n5), .ZN(n72) );
  AOI22_X1 U8 ( .A1(N127), .A2(net132681), .B1(N63), .B2(n5), .ZN(n73) );
  AOI22_X1 U9 ( .A1(N126), .A2(net132687), .B1(N62), .B2(n5), .ZN(n74) );
  BUF_X1 U10 ( .A(n9), .Z(n6) );
  BUF_X1 U11 ( .A(n6), .Z(net132697) );
  BUF_X1 U12 ( .A(n6), .Z(net132695) );
  BUF_X1 U13 ( .A(MUL_SGN_usgn), .Z(n9) );
  BUF_X1 U14 ( .A(n9), .Z(net132731) );
  BUF_X1 U15 ( .A(n9), .Z(net132729) );
  BUF_X1 U16 ( .A(n7), .Z(net132725) );
  BUF_X1 U17 ( .A(n8), .Z(n7) );
  BUF_X1 U18 ( .A(n7), .Z(net132723) );
  BUF_X1 U19 ( .A(MUL_SGN_usgn), .Z(n8) );
  BUF_X1 U20 ( .A(n8), .Z(net132735) );
  BUF_X1 U21 ( .A(n8), .Z(net132733) );
  INV_X1 U22 ( .A(net132725), .ZN(net132681) );
  INV_X1 U23 ( .A(net132725), .ZN(net132687) );
  INV_X1 U24 ( .A(net132725), .ZN(net132689) );
  BUF_X1 U25 ( .A(net132735), .Z(net132721) );
  BUF_X1 U26 ( .A(net132735), .Z(net132719) );
  BUF_X1 U27 ( .A(net132735), .Z(net132717) );
  BUF_X1 U28 ( .A(net132733), .Z(net132715) );
  BUF_X1 U29 ( .A(net132733), .Z(net132713) );
  BUF_X1 U30 ( .A(net132733), .Z(net132711) );
  BUF_X1 U31 ( .A(net132731), .Z(net132709) );
  BUF_X1 U32 ( .A(net132731), .Z(net132707) );
  BUF_X1 U33 ( .A(net132731), .Z(net132705) );
  BUF_X1 U34 ( .A(net132729), .Z(net132703) );
  BUF_X1 U35 ( .A(net132729), .Z(net132701) );
  BUF_X1 U36 ( .A(net132729), .Z(net132699) );
  INV_X1 U37 ( .A(n72), .ZN(N192) );
  INV_X1 U38 ( .A(n73), .ZN(N191) );
  INV_X1 U39 ( .A(n74), .ZN(N190) );
  INV_X1 U40 ( .A(n75), .ZN(N189) );
  AOI22_X1 U41 ( .A1(N125), .A2(net132689), .B1(N61), .B2(net132695), .ZN(n75)
         );
  INV_X1 U42 ( .A(n76), .ZN(N188) );
  AOI22_X1 U43 ( .A1(N124), .A2(net132689), .B1(N60), .B2(net132695), .ZN(n76)
         );
  INV_X1 U44 ( .A(n77), .ZN(N187) );
  AOI22_X1 U45 ( .A1(N123), .A2(net132689), .B1(N59), .B2(net132695), .ZN(n77)
         );
  INV_X1 U46 ( .A(n78), .ZN(N186) );
  AOI22_X1 U47 ( .A1(N122), .A2(net132689), .B1(N58), .B2(net132695), .ZN(n78)
         );
  INV_X1 U48 ( .A(n79), .ZN(N185) );
  AOI22_X1 U49 ( .A1(N121), .A2(net132689), .B1(N57), .B2(net132697), .ZN(n79)
         );
  INV_X1 U50 ( .A(n80), .ZN(N184) );
  AOI22_X1 U51 ( .A1(N120), .A2(net132689), .B1(N56), .B2(net132697), .ZN(n80)
         );
  INV_X1 U52 ( .A(n81), .ZN(N183) );
  AOI22_X1 U53 ( .A1(N119), .A2(net132689), .B1(N55), .B2(net132697), .ZN(n81)
         );
  INV_X1 U54 ( .A(n101), .ZN(N163) );
  AOI22_X1 U55 ( .A1(N99), .A2(net132681), .B1(N35), .B2(net132707), .ZN(n101)
         );
  INV_X1 U56 ( .A(n102), .ZN(N162) );
  AOI22_X1 U57 ( .A1(N98), .A2(net132689), .B1(N34), .B2(net132707), .ZN(n102)
         );
  INV_X1 U58 ( .A(n105), .ZN(N159) );
  AOI22_X1 U59 ( .A1(N95), .A2(net132689), .B1(N31), .B2(net132709), .ZN(n105)
         );
  INV_X1 U60 ( .A(n104), .ZN(N160) );
  AOI22_X1 U61 ( .A1(N96), .A2(net132681), .B1(N32), .B2(net132709), .ZN(n104)
         );
  INV_X1 U62 ( .A(n109), .ZN(N155) );
  AOI22_X1 U63 ( .A1(N91), .A2(net132687), .B1(N27), .B2(net132711), .ZN(n109)
         );
  INV_X1 U64 ( .A(n108), .ZN(N156) );
  AOI22_X1 U65 ( .A1(N92), .A2(net132689), .B1(N28), .B2(net132711), .ZN(n108)
         );
  INV_X1 U66 ( .A(n107), .ZN(N157) );
  AOI22_X1 U67 ( .A1(N93), .A2(net132681), .B1(N29), .B2(net132711), .ZN(n107)
         );
  INV_X1 U68 ( .A(n106), .ZN(N158) );
  AOI22_X1 U69 ( .A1(N94), .A2(net132687), .B1(N30), .B2(net132709), .ZN(n106)
         );
  INV_X1 U70 ( .A(n96), .ZN(N168) );
  AOI22_X1 U71 ( .A1(N104), .A2(net132687), .B1(N40), .B2(net132705), .ZN(n96)
         );
  INV_X1 U72 ( .A(n89), .ZN(N175) );
  AOI22_X1 U73 ( .A1(N111), .A2(net132687), .B1(N47), .B2(net132701), .ZN(n89)
         );
  INV_X1 U74 ( .A(n90), .ZN(N174) );
  AOI22_X1 U75 ( .A1(N110), .A2(net132687), .B1(N46), .B2(net132701), .ZN(n90)
         );
  INV_X1 U76 ( .A(n93), .ZN(N171) );
  AOI22_X1 U77 ( .A1(N107), .A2(net132687), .B1(N43), .B2(net132703), .ZN(n93)
         );
  INV_X1 U78 ( .A(n91), .ZN(N173) );
  AOI22_X1 U79 ( .A1(N109), .A2(net132687), .B1(N45), .B2(net132703), .ZN(n91)
         );
  INV_X1 U80 ( .A(n94), .ZN(N170) );
  AOI22_X1 U81 ( .A1(N106), .A2(net132687), .B1(N42), .B2(net132703), .ZN(n94)
         );
  INV_X1 U82 ( .A(n92), .ZN(N172) );
  AOI22_X1 U83 ( .A1(N108), .A2(net132687), .B1(N44), .B2(net132703), .ZN(n92)
         );
  INV_X1 U84 ( .A(n95), .ZN(N169) );
  AOI22_X1 U85 ( .A1(N105), .A2(net132687), .B1(N41), .B2(net132705), .ZN(n95)
         );
  INV_X1 U86 ( .A(n97), .ZN(N167) );
  AOI22_X1 U87 ( .A1(N103), .A2(net132687), .B1(N39), .B2(net132705), .ZN(n97)
         );
  INV_X1 U88 ( .A(n98), .ZN(N166) );
  AOI22_X1 U89 ( .A1(N102), .A2(net132687), .B1(N38), .B2(net132705), .ZN(n98)
         );
  INV_X1 U90 ( .A(n99), .ZN(N165) );
  AOI22_X1 U91 ( .A1(N101), .A2(net132689), .B1(N37), .B2(net132707), .ZN(n99)
         );
  INV_X1 U92 ( .A(n100), .ZN(N164) );
  AOI22_X1 U93 ( .A1(N100), .A2(net132687), .B1(N36), .B2(net132707), .ZN(n100) );
  INV_X1 U94 ( .A(n103), .ZN(N161) );
  AOI22_X1 U95 ( .A1(N97), .A2(net132689), .B1(N33), .B2(net132709), .ZN(n103)
         );
  INV_X1 U96 ( .A(n111), .ZN(N153) );
  AOI22_X1 U97 ( .A1(N89), .A2(net132687), .B1(N25), .B2(net132713), .ZN(n111)
         );
  INV_X1 U98 ( .A(n110), .ZN(N154) );
  AOI22_X1 U99 ( .A1(N90), .A2(net132687), .B1(N26), .B2(net132711), .ZN(n110)
         );
  INV_X1 U100 ( .A(n82), .ZN(N182) );
  AOI22_X1 U101 ( .A1(N118), .A2(net132689), .B1(N54), .B2(net132697), .ZN(n82) );
  INV_X1 U102 ( .A(n83), .ZN(N181) );
  AOI22_X1 U103 ( .A1(N117), .A2(net132689), .B1(N53), .B2(net132699), .ZN(n83) );
  INV_X1 U104 ( .A(n85), .ZN(N179) );
  AOI22_X1 U105 ( .A1(N115), .A2(net132689), .B1(N51), .B2(net132699), .ZN(n85) );
  INV_X1 U106 ( .A(n84), .ZN(N180) );
  AOI22_X1 U107 ( .A1(N116), .A2(net132689), .B1(N52), .B2(net132699), .ZN(n84) );
  INV_X1 U108 ( .A(n86), .ZN(N178) );
  AOI22_X1 U109 ( .A1(N114), .A2(net132689), .B1(N50), .B2(net132699), .ZN(n86) );
  INV_X1 U110 ( .A(n87), .ZN(N177) );
  AOI22_X1 U111 ( .A1(N113), .A2(net132687), .B1(N49), .B2(net132701), .ZN(n87) );
  INV_X1 U112 ( .A(n88), .ZN(N176) );
  AOI22_X1 U113 ( .A1(N112), .A2(net132687), .B1(N48), .B2(net132701), .ZN(n88) );
  INV_X1 U114 ( .A(n112), .ZN(N152) );
  AOI22_X1 U115 ( .A1(N88), .A2(net132681), .B1(N24), .B2(net132713), .ZN(n112) );
  INV_X1 U116 ( .A(n120), .ZN(N144) );
  AOI22_X1 U117 ( .A1(N80), .A2(net132689), .B1(N16), .B2(net132717), .ZN(n120) );
  INV_X1 U118 ( .A(n119), .ZN(N145) );
  AOI22_X1 U119 ( .A1(N81), .A2(net132681), .B1(N17), .B2(net132717), .ZN(n119) );
  INV_X1 U120 ( .A(n117), .ZN(N147) );
  AOI22_X1 U121 ( .A1(N83), .A2(net132687), .B1(N19), .B2(net132715), .ZN(n117) );
  INV_X1 U122 ( .A(n115), .ZN(N149) );
  AOI22_X1 U123 ( .A1(N85), .A2(net132681), .B1(N21), .B2(net132715), .ZN(n115) );
  INV_X1 U124 ( .A(n113), .ZN(N151) );
  AOI22_X1 U125 ( .A1(N87), .A2(net132689), .B1(N23), .B2(net132713), .ZN(n113) );
  INV_X1 U126 ( .A(n118), .ZN(N146) );
  AOI22_X1 U127 ( .A1(N82), .A2(net132681), .B1(N18), .B2(net132715), .ZN(n118) );
  INV_X1 U128 ( .A(n116), .ZN(N148) );
  AOI22_X1 U129 ( .A1(N84), .A2(net132687), .B1(N20), .B2(net132715), .ZN(n116) );
  INV_X1 U130 ( .A(n114), .ZN(N150) );
  AOI22_X1 U131 ( .A1(N86), .A2(net132687), .B1(N22), .B2(net132713), .ZN(n114) );
  INV_X1 U132 ( .A(n127), .ZN(N137) );
  AOI22_X1 U133 ( .A1(N73), .A2(net132681), .B1(N9), .B2(net132721), .ZN(n127)
         );
  INV_X1 U134 ( .A(n125), .ZN(N139) );
  AOI22_X1 U135 ( .A1(N75), .A2(net132681), .B1(N11), .B2(net132719), .ZN(n125) );
  INV_X1 U136 ( .A(n124), .ZN(N140) );
  AOI22_X1 U137 ( .A1(N76), .A2(net132681), .B1(N12), .B2(net132719), .ZN(n124) );
  INV_X1 U138 ( .A(n123), .ZN(N141) );
  AOI22_X1 U139 ( .A1(N77), .A2(net132681), .B1(N13), .B2(net132719), .ZN(n123) );
  INV_X1 U140 ( .A(n121), .ZN(N143) );
  AOI22_X1 U141 ( .A1(N79), .A2(net132689), .B1(N15), .B2(net132717), .ZN(n121) );
  INV_X1 U142 ( .A(n128), .ZN(N136) );
  AOI22_X1 U143 ( .A1(N72), .A2(net132681), .B1(N8), .B2(net132721), .ZN(n128)
         );
  INV_X1 U144 ( .A(n126), .ZN(N138) );
  AOI22_X1 U145 ( .A1(N74), .A2(net132681), .B1(N10), .B2(net132719), .ZN(n126) );
  INV_X1 U146 ( .A(n122), .ZN(N142) );
  AOI22_X1 U147 ( .A1(N78), .A2(net132681), .B1(N14), .B2(net132717), .ZN(n122) );
  INV_X1 U148 ( .A(n132), .ZN(N132) );
  AOI22_X1 U149 ( .A1(N68), .A2(net132681), .B1(N4), .B2(net132723), .ZN(n132)
         );
  INV_X1 U150 ( .A(n131), .ZN(N133) );
  AOI22_X1 U151 ( .A1(N69), .A2(net132681), .B1(N5), .B2(net132723), .ZN(n131)
         );
  INV_X1 U152 ( .A(n130), .ZN(N134) );
  AOI22_X1 U153 ( .A1(N70), .A2(net132681), .B1(N6), .B2(net132721), .ZN(n130)
         );
  INV_X1 U154 ( .A(n134), .ZN(N130) );
  AOI22_X1 U155 ( .A1(N66), .A2(net132681), .B1(N2), .B2(net132723), .ZN(n134)
         );
  INV_X1 U156 ( .A(n133), .ZN(N131) );
  AOI22_X1 U157 ( .A1(N67), .A2(net132681), .B1(N3), .B2(net132723), .ZN(n133)
         );
  INV_X1 U158 ( .A(n129), .ZN(N135) );
  AOI22_X1 U159 ( .A1(N71), .A2(net132681), .B1(N7), .B2(net132721), .ZN(n129)
         );
endmodule


module ALU_NBIT_ALU32_NBIT_BS_AMOUNT5 ( ALU_OpA, ALU_OpB, ALU_Opcode, 
        ALU_BS_amount, ALU_output, ALU_flags );
  input [31:0] ALU_OpA;
  input [31:0] ALU_OpB;
  input [5:0] ALU_Opcode;
  input [4:0] ALU_BS_amount;
  output [31:0] ALU_output;
  output [4:0] ALU_flags;
  wire   n19, s_P4_cin, s_from_P4_c_out, \s_mux_signals[1][0][31] ,
         \s_mux_signals[1][0][30] , \s_mux_signals[1][0][29] ,
         \s_mux_signals[1][0][28] , \s_mux_signals[1][0][27] ,
         \s_mux_signals[1][0][26] , \s_mux_signals[1][0][25] ,
         \s_mux_signals[1][0][24] , \s_mux_signals[1][0][23] ,
         \s_mux_signals[1][0][22] , \s_mux_signals[1][0][21] ,
         \s_mux_signals[1][0][20] , \s_mux_signals[1][0][19] ,
         \s_mux_signals[1][0][18] , \s_mux_signals[1][0][17] ,
         \s_mux_signals[1][0][16] , \s_mux_signals[1][0][15] ,
         \s_mux_signals[1][0][14] , \s_mux_signals[1][0][13] ,
         \s_mux_signals[1][0][12] , \s_mux_signals[1][0][11] ,
         \s_mux_signals[1][0][10] , \s_mux_signals[1][0][9] ,
         \s_mux_signals[1][0][8] , \s_mux_signals[1][0][7] ,
         \s_mux_signals[1][0][6] , \s_mux_signals[1][0][5] ,
         \s_mux_signals[1][0][4] , \s_mux_signals[1][0][3] ,
         \s_mux_signals[1][0][2] , \s_mux_signals[1][0][1] ,
         \s_mux_signals[1][0][0] , \s_mux_signals[1][1][31] ,
         \s_mux_signals[1][1][30] , \s_mux_signals[1][1][29] ,
         \s_mux_signals[1][1][28] , \s_mux_signals[1][1][27] ,
         \s_mux_signals[1][1][26] , \s_mux_signals[1][1][25] ,
         \s_mux_signals[1][1][24] , \s_mux_signals[1][1][23] ,
         \s_mux_signals[1][1][22] , \s_mux_signals[1][1][21] ,
         \s_mux_signals[1][1][20] , \s_mux_signals[1][1][19] ,
         \s_mux_signals[1][1][18] , \s_mux_signals[1][1][17] ,
         \s_mux_signals[1][1][16] , \s_mux_signals[1][1][15] ,
         \s_mux_signals[1][1][14] , \s_mux_signals[1][1][13] ,
         \s_mux_signals[1][1][12] , \s_mux_signals[1][1][11] ,
         \s_mux_signals[1][1][10] , \s_mux_signals[1][1][9] ,
         \s_mux_signals[1][1][8] , \s_mux_signals[1][1][7] ,
         \s_mux_signals[1][1][6] , \s_mux_signals[1][1][5] ,
         \s_mux_signals[1][1][4] , \s_mux_signals[1][1][3] ,
         \s_mux_signals[1][1][2] , \s_mux_signals[1][1][1] ,
         \s_mux_signals[1][1][0] , s_SGN_usgn, n39, n41, n42, n43, n44, n45,
         n46, n48, n11, n12, n14, n15, n16, n17, n18;
  wire   [1:0] s_BS_opcode;
  wire   [31:0] s_from_BS_to_units_opA;
  wire   [31:0] s_OpB;
  wire   [31:0] s_not_opB;
  wire   [31:0] s_sel_opB;
  wire   [31:0] s_from_P4_to_out_sum;
  wire   [3:0] s_LU_opcode;
  wire   [31:0] s_from_LU_to_out_mux;
  wire   [3:0] s_CMP_opcode;
  wire   [31:0] s_from_CMP_to_out_mux;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30;

  NOR2_X2 U83 ( .A1(n44), .A2(n39), .ZN(s_BS_opcode[1]) );
  OR2_X2 U86 ( .A1(ALU_Opcode[4]), .A2(ALU_Opcode[5]), .ZN(n39) );
  Barrel_Shifter_NBIT_AMOUNT5 BS ( .BS_data_in(ALU_OpA), .BS_opcode(
        s_BS_opcode), .BS_amount(ALU_BS_amount), .BS_data_out(
        s_from_BS_to_units_opA) );
  Mux_NBit_2x1_NBIT_IN32_15 MuxP4 ( .port0(s_OpB), .port1(s_not_opB), .sel(
        s_P4_cin), .portY(s_sel_opB) );
  P4Adder_N32 P4 ( .A({n12, n11, s_from_BS_to_units_opA[29:0]}), .B(s_sel_opB), 
        .c_in(s_P4_cin), .c_out(s_from_P4_c_out), .Sum(s_from_P4_to_out_sum)
         );
  Logic_Unit_NBIT_DATA32 LU ( .LU_OpA({n12, n11, s_from_BS_to_units_opA[29:0]}), .LU_OpB(ALU_OpB), .LU_Opcode(s_LU_opcode), .LU_Y(s_from_LU_to_out_mux) );
  Comparison_Logic_NBIT_DATA32 CMPL ( .CMPL_OpA(s_from_BS_to_units_opA), 
        .CMPL_OpB(ALU_OpB), .CMPL_OPCODE(s_CMP_opcode), .CMPL_Y({
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15, 
        SYNOPSYS_UNCONNECTED__16, SYNOPSYS_UNCONNECTED__17, 
        SYNOPSYS_UNCONNECTED__18, SYNOPSYS_UNCONNECTED__19, 
        SYNOPSYS_UNCONNECTED__20, SYNOPSYS_UNCONNECTED__21, 
        SYNOPSYS_UNCONNECTED__22, SYNOPSYS_UNCONNECTED__23, 
        SYNOPSYS_UNCONNECTED__24, SYNOPSYS_UNCONNECTED__25, 
        SYNOPSYS_UNCONNECTED__26, SYNOPSYS_UNCONNECTED__27, 
        SYNOPSYS_UNCONNECTED__28, SYNOPSYS_UNCONNECTED__29, 
        SYNOPSYS_UNCONNECTED__30, s_from_CMP_to_out_mux[0]}) );
  Mux_NBit_2x1_NBIT_IN32_14 MUX1 ( .port0(s_from_P4_to_out_sum), .port1(
        s_from_LU_to_out_mux), .sel(ALU_Opcode[4]), .portY({
        \s_mux_signals[1][0][31] , \s_mux_signals[1][0][30] , 
        \s_mux_signals[1][0][29] , \s_mux_signals[1][0][28] , 
        \s_mux_signals[1][0][27] , \s_mux_signals[1][0][26] , 
        \s_mux_signals[1][0][25] , \s_mux_signals[1][0][24] , 
        \s_mux_signals[1][0][23] , \s_mux_signals[1][0][22] , 
        \s_mux_signals[1][0][21] , \s_mux_signals[1][0][20] , 
        \s_mux_signals[1][0][19] , \s_mux_signals[1][0][18] , 
        \s_mux_signals[1][0][17] , \s_mux_signals[1][0][16] , 
        \s_mux_signals[1][0][15] , \s_mux_signals[1][0][14] , 
        \s_mux_signals[1][0][13] , \s_mux_signals[1][0][12] , 
        \s_mux_signals[1][0][11] , \s_mux_signals[1][0][10] , 
        \s_mux_signals[1][0][9] , \s_mux_signals[1][0][8] , 
        \s_mux_signals[1][0][7] , \s_mux_signals[1][0][6] , 
        \s_mux_signals[1][0][5] , \s_mux_signals[1][0][4] , 
        \s_mux_signals[1][0][3] , \s_mux_signals[1][0][2] , 
        \s_mux_signals[1][0][1] , \s_mux_signals[1][0][0] }) );
  Mux_NBit_2x1_NBIT_IN32_13 MUX2 ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, s_from_CMP_to_out_mux[0]}), .port1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .sel(ALU_Opcode[4]), .portY({
        \s_mux_signals[1][1][31] , \s_mux_signals[1][1][30] , 
        \s_mux_signals[1][1][29] , \s_mux_signals[1][1][28] , 
        \s_mux_signals[1][1][27] , \s_mux_signals[1][1][26] , 
        \s_mux_signals[1][1][25] , \s_mux_signals[1][1][24] , 
        \s_mux_signals[1][1][23] , \s_mux_signals[1][1][22] , 
        \s_mux_signals[1][1][21] , \s_mux_signals[1][1][20] , 
        \s_mux_signals[1][1][19] , \s_mux_signals[1][1][18] , 
        \s_mux_signals[1][1][17] , \s_mux_signals[1][1][16] , 
        \s_mux_signals[1][1][15] , \s_mux_signals[1][1][14] , 
        \s_mux_signals[1][1][13] , \s_mux_signals[1][1][12] , 
        \s_mux_signals[1][1][11] , \s_mux_signals[1][1][10] , 
        \s_mux_signals[1][1][9] , \s_mux_signals[1][1][8] , 
        \s_mux_signals[1][1][7] , \s_mux_signals[1][1][6] , 
        \s_mux_signals[1][1][5] , \s_mux_signals[1][1][4] , 
        \s_mux_signals[1][1][3] , \s_mux_signals[1][1][2] , 
        \s_mux_signals[1][1][1] , \s_mux_signals[1][1][0] }) );
  Mux_NBit_2x1_NBIT_IN32_12 MUX3 ( .port0({\s_mux_signals[1][0][31] , 
        \s_mux_signals[1][0][30] , \s_mux_signals[1][0][29] , 
        \s_mux_signals[1][0][28] , \s_mux_signals[1][0][27] , 
        \s_mux_signals[1][0][26] , \s_mux_signals[1][0][25] , 
        \s_mux_signals[1][0][24] , \s_mux_signals[1][0][23] , 
        \s_mux_signals[1][0][22] , \s_mux_signals[1][0][21] , 
        \s_mux_signals[1][0][20] , \s_mux_signals[1][0][19] , 
        \s_mux_signals[1][0][18] , \s_mux_signals[1][0][17] , 
        \s_mux_signals[1][0][16] , \s_mux_signals[1][0][15] , 
        \s_mux_signals[1][0][14] , \s_mux_signals[1][0][13] , 
        \s_mux_signals[1][0][12] , \s_mux_signals[1][0][11] , 
        \s_mux_signals[1][0][10] , \s_mux_signals[1][0][9] , 
        \s_mux_signals[1][0][8] , \s_mux_signals[1][0][7] , 
        \s_mux_signals[1][0][6] , \s_mux_signals[1][0][5] , 
        \s_mux_signals[1][0][4] , \s_mux_signals[1][0][3] , 
        \s_mux_signals[1][0][2] , \s_mux_signals[1][0][1] , 
        \s_mux_signals[1][0][0] }), .port1({\s_mux_signals[1][1][31] , 
        \s_mux_signals[1][1][30] , \s_mux_signals[1][1][29] , 
        \s_mux_signals[1][1][28] , \s_mux_signals[1][1][27] , 
        \s_mux_signals[1][1][26] , \s_mux_signals[1][1][25] , 
        \s_mux_signals[1][1][24] , \s_mux_signals[1][1][23] , 
        \s_mux_signals[1][1][22] , \s_mux_signals[1][1][21] , 
        \s_mux_signals[1][1][20] , \s_mux_signals[1][1][19] , 
        \s_mux_signals[1][1][18] , \s_mux_signals[1][1][17] , 
        \s_mux_signals[1][1][16] , \s_mux_signals[1][1][15] , 
        \s_mux_signals[1][1][14] , \s_mux_signals[1][1][13] , 
        \s_mux_signals[1][1][12] , \s_mux_signals[1][1][11] , 
        \s_mux_signals[1][1][10] , \s_mux_signals[1][1][9] , 
        \s_mux_signals[1][1][8] , \s_mux_signals[1][1][7] , 
        \s_mux_signals[1][1][6] , \s_mux_signals[1][1][5] , 
        \s_mux_signals[1][1][4] , \s_mux_signals[1][1][3] , 
        \s_mux_signals[1][1][2] , \s_mux_signals[1][1][1] , 
        \s_mux_signals[1][1][0] }), .sel(ALU_Opcode[5]), .portY({
        ALU_output[31:1], n19}) );
  Flag_Generator_NBIT_ALU32 FG ( .FG_ALU_out({ALU_output[31:1], n19}), 
        .FG_sgn_usgn(s_SGN_usgn), .FG_carry(s_from_P4_c_out), .FG_ZF(
        ALU_flags[0]), .FG_PF(ALU_flags[1]), .FG_SF(ALU_flags[2]), .FG_CF(
        ALU_flags[3]), .FG_OF(ALU_flags[4]) );
  NOR2_X1 U2 ( .A1(n39), .A2(n42), .ZN(s_P4_cin) );
  CLKBUF_X1 U3 ( .A(s_from_BS_to_units_opA[30]), .Z(n11) );
  BUF_X1 U4 ( .A(n43), .Z(n14) );
  BUF_X1 U5 ( .A(n43), .Z(n15) );
  BUF_X1 U6 ( .A(n43), .Z(n16) );
  INV_X1 U7 ( .A(s_not_opB[6]), .ZN(s_OpB[6]) );
  NAND2_X1 U8 ( .A1(ALU_OpB[6]), .A2(n16), .ZN(s_not_opB[6]) );
  INV_X1 U9 ( .A(s_not_opB[2]), .ZN(s_OpB[2]) );
  NAND2_X1 U10 ( .A1(ALU_OpB[2]), .A2(n15), .ZN(s_not_opB[2]) );
  INV_X1 U11 ( .A(s_not_opB[4]), .ZN(s_OpB[4]) );
  NAND2_X1 U12 ( .A1(ALU_OpB[4]), .A2(n16), .ZN(s_not_opB[4]) );
  INV_X1 U13 ( .A(s_not_opB[5]), .ZN(s_OpB[5]) );
  NAND2_X1 U14 ( .A1(ALU_OpB[5]), .A2(n16), .ZN(s_not_opB[5]) );
  INV_X1 U15 ( .A(s_not_opB[3]), .ZN(s_OpB[3]) );
  NAND2_X1 U16 ( .A1(ALU_OpB[3]), .A2(n16), .ZN(s_not_opB[3]) );
  INV_X1 U17 ( .A(s_not_opB[7]), .ZN(s_OpB[7]) );
  NAND2_X1 U18 ( .A1(ALU_OpB[7]), .A2(n16), .ZN(s_not_opB[7]) );
  INV_X1 U19 ( .A(s_not_opB[9]), .ZN(s_OpB[9]) );
  NAND2_X1 U20 ( .A1(ALU_OpB[9]), .A2(n16), .ZN(s_not_opB[9]) );
  INV_X1 U21 ( .A(s_not_opB[17]), .ZN(s_OpB[17]) );
  NAND2_X1 U22 ( .A1(ALU_OpB[17]), .A2(n14), .ZN(s_not_opB[17]) );
  INV_X1 U23 ( .A(s_not_opB[16]), .ZN(s_OpB[16]) );
  NAND2_X1 U24 ( .A1(ALU_OpB[16]), .A2(n14), .ZN(s_not_opB[16]) );
  INV_X1 U25 ( .A(s_not_opB[0]), .ZN(s_OpB[0]) );
  NAND2_X1 U26 ( .A1(ALU_OpB[0]), .A2(n14), .ZN(s_not_opB[0]) );
  INV_X1 U27 ( .A(s_not_opB[13]), .ZN(s_OpB[13]) );
  NAND2_X1 U28 ( .A1(ALU_OpB[13]), .A2(n14), .ZN(s_not_opB[13]) );
  INV_X1 U29 ( .A(s_not_opB[25]), .ZN(s_OpB[25]) );
  NAND2_X1 U30 ( .A1(ALU_OpB[25]), .A2(n15), .ZN(s_not_opB[25]) );
  INV_X1 U31 ( .A(s_not_opB[12]), .ZN(s_OpB[12]) );
  NAND2_X1 U32 ( .A1(ALU_OpB[12]), .A2(n14), .ZN(s_not_opB[12]) );
  INV_X1 U33 ( .A(s_not_opB[10]), .ZN(s_OpB[10]) );
  NAND2_X1 U34 ( .A1(ALU_OpB[10]), .A2(n14), .ZN(s_not_opB[10]) );
  INV_X1 U35 ( .A(s_not_opB[20]), .ZN(s_OpB[20]) );
  NAND2_X1 U36 ( .A1(ALU_OpB[20]), .A2(n15), .ZN(s_not_opB[20]) );
  INV_X1 U37 ( .A(s_not_opB[21]), .ZN(s_OpB[21]) );
  NAND2_X1 U38 ( .A1(ALU_OpB[21]), .A2(n15), .ZN(s_not_opB[21]) );
  INV_X1 U39 ( .A(s_not_opB[22]), .ZN(s_OpB[22]) );
  NAND2_X1 U40 ( .A1(ALU_OpB[22]), .A2(n15), .ZN(s_not_opB[22]) );
  INV_X1 U41 ( .A(s_not_opB[18]), .ZN(s_OpB[18]) );
  NAND2_X1 U42 ( .A1(ALU_OpB[18]), .A2(n14), .ZN(s_not_opB[18]) );
  INV_X1 U43 ( .A(s_not_opB[1]), .ZN(s_OpB[1]) );
  NAND2_X1 U44 ( .A1(ALU_OpB[1]), .A2(n14), .ZN(s_not_opB[1]) );
  INV_X1 U45 ( .A(s_not_opB[14]), .ZN(s_OpB[14]) );
  NAND2_X1 U46 ( .A1(ALU_OpB[14]), .A2(n14), .ZN(s_not_opB[14]) );
  INV_X1 U47 ( .A(s_not_opB[28]), .ZN(s_OpB[28]) );
  NAND2_X1 U48 ( .A1(ALU_OpB[28]), .A2(n15), .ZN(s_not_opB[28]) );
  INV_X1 U49 ( .A(s_not_opB[29]), .ZN(s_OpB[29]) );
  NAND2_X1 U50 ( .A1(ALU_OpB[29]), .A2(n15), .ZN(s_not_opB[29]) );
  INV_X1 U51 ( .A(s_not_opB[24]), .ZN(s_OpB[24]) );
  NAND2_X1 U52 ( .A1(ALU_OpB[24]), .A2(n15), .ZN(s_not_opB[24]) );
  INV_X1 U53 ( .A(s_not_opB[26]), .ZN(s_OpB[26]) );
  NAND2_X1 U54 ( .A1(ALU_OpB[26]), .A2(n15), .ZN(s_not_opB[26]) );
  INV_X1 U55 ( .A(s_not_opB[8]), .ZN(s_OpB[8]) );
  NAND2_X1 U56 ( .A1(ALU_OpB[8]), .A2(n16), .ZN(s_not_opB[8]) );
  INV_X1 U57 ( .A(s_not_opB[11]), .ZN(s_OpB[11]) );
  NAND2_X1 U58 ( .A1(ALU_OpB[11]), .A2(n14), .ZN(s_not_opB[11]) );
  INV_X1 U59 ( .A(s_not_opB[15]), .ZN(s_OpB[15]) );
  NAND2_X1 U60 ( .A1(ALU_OpB[15]), .A2(n14), .ZN(s_not_opB[15]) );
  INV_X1 U61 ( .A(s_not_opB[19]), .ZN(s_OpB[19]) );
  NAND2_X1 U62 ( .A1(ALU_OpB[19]), .A2(n14), .ZN(s_not_opB[19]) );
  INV_X1 U63 ( .A(s_not_opB[23]), .ZN(s_OpB[23]) );
  NAND2_X1 U64 ( .A1(ALU_OpB[23]), .A2(n15), .ZN(s_not_opB[23]) );
  INV_X1 U65 ( .A(s_not_opB[27]), .ZN(s_OpB[27]) );
  NAND2_X1 U66 ( .A1(ALU_OpB[27]), .A2(n15), .ZN(s_not_opB[27]) );
  INV_X1 U67 ( .A(s_not_opB[30]), .ZN(s_OpB[30]) );
  NAND2_X1 U68 ( .A1(ALU_OpB[30]), .A2(n15), .ZN(s_not_opB[30]) );
  INV_X1 U69 ( .A(s_not_opB[31]), .ZN(s_OpB[31]) );
  NAND2_X1 U70 ( .A1(ALU_OpB[31]), .A2(n16), .ZN(s_not_opB[31]) );
  NOR2_X1 U71 ( .A1(s_BS_opcode[0]), .A2(s_BS_opcode[1]), .ZN(n43) );
  NOR2_X1 U72 ( .A1(n17), .A2(n48), .ZN(s_CMP_opcode[1]) );
  NOR2_X1 U73 ( .A1(n17), .A2(n45), .ZN(s_LU_opcode[1]) );
  OAI21_X1 U74 ( .B1(n39), .B2(n17), .A(n41), .ZN(s_SGN_usgn) );
  INV_X1 U75 ( .A(s_CMP_opcode[3]), .ZN(n41) );
  NOR2_X1 U76 ( .A1(n46), .A2(n39), .ZN(s_BS_opcode[0]) );
  NOR2_X1 U77 ( .A1(n48), .A2(n42), .ZN(s_CMP_opcode[0]) );
  NOR2_X1 U78 ( .A1(n46), .A2(n45), .ZN(s_LU_opcode[2]) );
  NOR2_X1 U79 ( .A1(n44), .A2(n45), .ZN(s_LU_opcode[3]) );
  NAND2_X1 U80 ( .A1(ALU_Opcode[4]), .A2(n18), .ZN(n45) );
  NOR2_X1 U81 ( .A1(n46), .A2(n48), .ZN(s_CMP_opcode[2]) );
  NOR2_X1 U82 ( .A1(n42), .A2(n45), .ZN(s_LU_opcode[0]) );
  OR2_X1 U84 ( .A1(n18), .A2(ALU_Opcode[4]), .ZN(n48) );
  NOR2_X1 U85 ( .A1(n48), .A2(n44), .ZN(s_CMP_opcode[3]) );
  INV_X1 U87 ( .A(ALU_Opcode[5]), .ZN(n18) );
  INV_X1 U119 ( .A(ALU_Opcode[3]), .ZN(n44) );
  INV_X1 U120 ( .A(ALU_Opcode[2]), .ZN(n46) );
  INV_X1 U121 ( .A(ALU_Opcode[0]), .ZN(n42) );
  CLKBUF_X1 U122 ( .A(s_from_BS_to_units_opA[31]), .Z(n12) );
  CLKBUF_X1 U123 ( .A(n19), .Z(ALU_output[0]) );
  INV_X1 U124 ( .A(ALU_Opcode[1]), .ZN(n17) );
endmodule


module Enable_Interface_NBIT_DATA32_0 ( EI_datain, EI_enable, EI_dataout );
  input [31:0] EI_datain;
  output [31:0] EI_dataout;
  input EI_enable;
  wire   n1, n2, n3;

  BUF_X1 U1 ( .A(EI_enable), .Z(n3) );
  BUF_X1 U2 ( .A(EI_enable), .Z(n2) );
  BUF_X1 U3 ( .A(EI_enable), .Z(n1) );
  AND2_X1 U4 ( .A1(EI_datain[17]), .A2(n1), .ZN(EI_dataout[17]) );
  AND2_X1 U5 ( .A1(EI_datain[18]), .A2(n1), .ZN(EI_dataout[18]) );
  AND2_X1 U6 ( .A1(EI_datain[19]), .A2(n1), .ZN(EI_dataout[19]) );
  AND2_X1 U7 ( .A1(EI_datain[16]), .A2(n1), .ZN(EI_dataout[16]) );
  AND2_X1 U8 ( .A1(EI_datain[21]), .A2(n2), .ZN(EI_dataout[21]) );
  AND2_X1 U9 ( .A1(EI_datain[20]), .A2(n2), .ZN(EI_dataout[20]) );
  AND2_X1 U10 ( .A1(EI_datain[23]), .A2(n2), .ZN(EI_dataout[23]) );
  AND2_X1 U11 ( .A1(EI_datain[24]), .A2(n2), .ZN(EI_dataout[24]) );
  AND2_X1 U12 ( .A1(EI_datain[26]), .A2(n2), .ZN(EI_dataout[26]) );
  AND2_X1 U13 ( .A1(EI_datain[25]), .A2(n2), .ZN(EI_dataout[25]) );
  AND2_X1 U14 ( .A1(EI_datain[27]), .A2(n2), .ZN(EI_dataout[27]) );
  AND2_X1 U15 ( .A1(EI_datain[28]), .A2(n2), .ZN(EI_dataout[28]) );
  AND2_X1 U16 ( .A1(EI_datain[29]), .A2(n2), .ZN(EI_dataout[29]) );
  AND2_X1 U17 ( .A1(EI_datain[15]), .A2(n1), .ZN(EI_dataout[15]) );
  AND2_X1 U18 ( .A1(EI_datain[0]), .A2(n1), .ZN(EI_dataout[0]) );
  AND2_X1 U19 ( .A1(EI_datain[2]), .A2(n2), .ZN(EI_dataout[2]) );
  AND2_X1 U20 ( .A1(EI_datain[1]), .A2(n1), .ZN(EI_dataout[1]) );
  AND2_X1 U21 ( .A1(EI_datain[5]), .A2(n3), .ZN(EI_dataout[5]) );
  AND2_X1 U22 ( .A1(EI_datain[4]), .A2(n3), .ZN(EI_dataout[4]) );
  AND2_X1 U23 ( .A1(EI_datain[3]), .A2(n3), .ZN(EI_dataout[3]) );
  AND2_X1 U24 ( .A1(EI_datain[13]), .A2(n1), .ZN(EI_dataout[13]) );
  AND2_X1 U25 ( .A1(EI_datain[10]), .A2(n1), .ZN(EI_dataout[10]) );
  AND2_X1 U26 ( .A1(EI_datain[11]), .A2(n1), .ZN(EI_dataout[11]) );
  AND2_X1 U27 ( .A1(EI_datain[12]), .A2(n1), .ZN(EI_dataout[12]) );
  AND2_X1 U28 ( .A1(EI_datain[14]), .A2(n1), .ZN(EI_dataout[14]) );
  AND2_X1 U29 ( .A1(n3), .A2(EI_datain[9]), .ZN(EI_dataout[9]) );
  AND2_X1 U30 ( .A1(EI_datain[8]), .A2(n3), .ZN(EI_dataout[8]) );
  AND2_X1 U31 ( .A1(EI_datain[22]), .A2(n2), .ZN(EI_dataout[22]) );
  AND2_X1 U32 ( .A1(EI_datain[7]), .A2(n3), .ZN(EI_dataout[7]) );
  AND2_X1 U33 ( .A1(EI_datain[6]), .A2(n3), .ZN(EI_dataout[6]) );
  AND2_X1 U34 ( .A1(EI_datain[30]), .A2(n2), .ZN(EI_dataout[30]) );
  AND2_X2 U35 ( .A1(EI_datain[31]), .A2(n3), .ZN(EI_dataout[31]) );
endmodule


module Jmp_Branch_Manager_N32 ( JBM_iszero, JBM_Reg, JBM_Imm, JBM_NPC, 
        JBM_JMP_branch, JBM_transparent_mode, JBM_Upd_PC, JBM_taken );
  input [31:0] JBM_Reg;
  input [31:0] JBM_Imm;
  input [31:0] JBM_NPC;
  input [1:0] JBM_JMP_branch;
  output [31:0] JBM_Upd_PC;
  input JBM_iszero, JBM_transparent_mode;
  output JBM_taken;
  wire   s_sel_muxes, n2, n3;
  wire   [31:0] s_Fmuxtrg_Tadd;
  wire   [31:0] s_Fmuxtba_Tadd;

  XOR2_X1 U5 ( .A(JBM_iszero), .B(JBM_JMP_branch[0]), .Z(n2) );
  Mux_NBit_2x1_NBIT_IN32_17 MUX_TRG ( .port0(JBM_Reg), .port1(JBM_Imm), .sel(
        s_sel_muxes), .portY(s_Fmuxtrg_Tadd) );
  Mux_NBit_2x1_NBIT_IN32_16 MUX_TBA ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .port1(JBM_NPC), .sel(s_sel_muxes), .portY(
        s_Fmuxtba_Tadd) );
  PropagateCarryLookahead_N32_1 ADD ( .A(s_Fmuxtrg_Tadd), .B(s_Fmuxtba_Tadd), 
        .Cin(1'b0), .Sum(JBM_Upd_PC) );
  OAI21_X1 U2 ( .B1(JBM_transparent_mode), .B2(n2), .A(n3), .ZN(JBM_taken) );
  INV_X1 U3 ( .A(JBM_JMP_branch[1]), .ZN(n3) );
  NAND2_X1 U4 ( .A1(JBM_JMP_branch[1]), .A2(JBM_JMP_branch[0]), .ZN(
        s_sel_muxes) );
endmodule


module NComparatorWithEnable_NBIT32_1 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13;

  ComparatorWithEnable_32 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n11), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_31 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n11), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_30 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n11), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_29 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n11), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_28 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n11), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_27 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n11), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_26 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n11), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_25 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n11), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_24 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n11), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_23 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n11), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_22 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n11), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_21 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n11), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_20 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n12), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_19 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n12), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_18 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n12), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_17 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n12), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_16 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n12), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_15 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n12), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_14 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n12), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_13 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n12), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_12 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n12), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_11 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n12), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_10 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n12), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_9 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n12), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_8 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n13), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_7 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n13), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_6 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n13), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_5 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n13), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_4 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n13), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_3 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n13), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_2 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n13), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_1 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n13), .y(
        \matrix[31][0] ) );
  NAND4_X1 U1 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n10) );
  NAND4_X1 U2 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n6) );
  NAND4_X1 U3 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n9) );
  NAND4_X1 U4 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(\matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n5) );
  NAND4_X1 U5 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(\matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n8) );
  NAND4_X1 U6 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n4) );
  NAND4_X1 U7 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n7) );
  AND2_X1 U8 ( .A1(n1), .A2(n2), .ZN(ComparatorBit) );
  NOR4_X1 U9 ( .A1(n3), .A2(n4), .A3(n5), .A4(n6), .ZN(n2) );
  NOR4_X1 U10 ( .A1(n7), .A2(n8), .A3(n9), .A4(n10), .ZN(n1) );
  NAND4_X1 U11 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n3) );
  CLKBUF_X1 U12 ( .A(Enable), .Z(n12) );
  CLKBUF_X1 U13 ( .A(Enable), .Z(n11) );
  CLKBUF_X1 U14 ( .A(Enable), .Z(n13) );
endmodule


module Sign_Extender_NBIT_DATA32 ( SE_I_J, SE_S_U, SE_in, SE_out );
  input [31:0] SE_in;
  output [31:0] SE_out;
  input SE_I_J, SE_S_U;
  wire   \SE_in[15] , \SE_in[14] , \SE_in[13] , \SE_in[12] , \SE_in[11] ,
         \SE_in[10] , \SE_in[9] , \SE_in[8] , \SE_in[7] , \SE_in[6] ,
         \SE_in[5] , \SE_in[4] , \SE_in[3] , \SE_in[2] , \SE_in[1] ,
         \SE_in[0] , s_and1, s_and2;
  wire   [25:16] s_tmp1;
  wire   [31:26] s_tmp2;
  assign SE_out[15] = \SE_in[15] ;
  assign \SE_in[15]  = SE_in[15];
  assign SE_out[14] = \SE_in[14] ;
  assign \SE_in[14]  = SE_in[14];
  assign SE_out[13] = \SE_in[13] ;
  assign \SE_in[13]  = SE_in[13];
  assign SE_out[12] = \SE_in[12] ;
  assign \SE_in[12]  = SE_in[12];
  assign SE_out[11] = \SE_in[11] ;
  assign \SE_in[11]  = SE_in[11];
  assign SE_out[10] = \SE_in[10] ;
  assign \SE_in[10]  = SE_in[10];
  assign SE_out[9] = \SE_in[9] ;
  assign \SE_in[9]  = SE_in[9];
  assign SE_out[8] = \SE_in[8] ;
  assign \SE_in[8]  = SE_in[8];
  assign SE_out[7] = \SE_in[7] ;
  assign \SE_in[7]  = SE_in[7];
  assign SE_out[6] = \SE_in[6] ;
  assign \SE_in[6]  = SE_in[6];
  assign SE_out[5] = \SE_in[5] ;
  assign \SE_in[5]  = SE_in[5];
  assign SE_out[4] = \SE_in[4] ;
  assign \SE_in[4]  = SE_in[4];
  assign SE_out[3] = \SE_in[3] ;
  assign \SE_in[3]  = SE_in[3];
  assign SE_out[2] = \SE_in[2] ;
  assign \SE_in[2]  = SE_in[2];
  assign SE_out[1] = \SE_in[1] ;
  assign \SE_in[1]  = SE_in[1];
  assign SE_out[0] = \SE_in[0] ;
  assign \SE_in[0]  = SE_in[0];

  Mux_NBit_2x1_NBIT_IN10_0 MUX_IMM ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .port1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .sel(s_and1), .portY(s_tmp1) );
  Mux_NBit_2x1_NBIT_IN6_0 MUX_JMP ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .port1({1'b1, 1'b1, 1'b1, 1'b1, 1'b1, 1'b1}), .sel(s_and2), .portY(s_tmp2)
         );
  Mux_NBit_2x1_NBIT_IN10_1 MUX_IMM_OUT ( .port0(SE_in[25:16]), .port1(s_tmp1), 
        .sel(SE_I_J), .portY(SE_out[25:16]) );
  Mux_NBit_2x1_NBIT_IN6_1 MUX_JMP_OUT ( .port0(s_tmp2), .port1(SE_out[25:20]), 
        .sel(SE_I_J), .portY(SE_out[31:26]) );
  AND2_X1 U3 ( .A1(\SE_in[15] ), .A2(SE_S_U), .ZN(s_and1) );
  AND2_X1 U4 ( .A1(SE_in[25]), .A2(SE_S_U), .ZN(s_and2) );
endmodule


module Register_File_NBIT_ADDR5_NBIT_DATA32 ( RF_clk, RF_reset, RF_enable, 
        RF_RD1, RF_RD2, RF_WR, RF_AddrRd1, RF_AddrRd2, RF_AddrWr, RF_data_in, 
        RF_out1, RF_out2 );
  input [4:0] RF_AddrRd1;
  input [4:0] RF_AddrRd2;
  input [4:0] RF_AddrWr;
  input [31:0] RF_data_in;
  output [31:0] RF_out1;
  output [31:0] RF_out2;
  input RF_clk, RF_reset, RF_enable, RF_RD1, RF_RD2, RF_WR;
  wire   s_wr_enable, s_rd1_enable, s_rd2_enable, \s_mux2_signals[0][0][31] ,
         \s_mux2_signals[0][0][30] , \s_mux2_signals[0][0][29] ,
         \s_mux2_signals[0][0][28] , \s_mux2_signals[0][0][27] ,
         \s_mux2_signals[0][0][26] , \s_mux2_signals[0][0][25] ,
         \s_mux2_signals[0][0][24] , \s_mux2_signals[0][0][23] ,
         \s_mux2_signals[0][0][22] , \s_mux2_signals[0][0][21] ,
         \s_mux2_signals[0][0][20] , \s_mux2_signals[0][0][19] ,
         \s_mux2_signals[0][0][18] , \s_mux2_signals[0][0][17] ,
         \s_mux2_signals[0][0][16] , \s_mux2_signals[0][0][15] ,
         \s_mux2_signals[0][0][14] , \s_mux2_signals[0][0][13] ,
         \s_mux2_signals[0][0][12] , \s_mux2_signals[0][0][11] ,
         \s_mux2_signals[0][0][10] , \s_mux2_signals[0][0][9] ,
         \s_mux2_signals[0][0][8] , \s_mux2_signals[0][0][7] ,
         \s_mux2_signals[0][0][6] , \s_mux2_signals[0][0][5] ,
         \s_mux2_signals[0][0][4] , \s_mux2_signals[0][0][3] ,
         \s_mux2_signals[0][0][2] , \s_mux2_signals[0][0][1] ,
         \s_mux2_signals[0][0][0] , \s_mux2_signals[0][1][31] ,
         \s_mux2_signals[0][1][30] , \s_mux2_signals[0][1][29] ,
         \s_mux2_signals[0][1][28] , \s_mux2_signals[0][1][27] ,
         \s_mux2_signals[0][1][26] , \s_mux2_signals[0][1][25] ,
         \s_mux2_signals[0][1][24] , \s_mux2_signals[0][1][23] ,
         \s_mux2_signals[0][1][22] , \s_mux2_signals[0][1][21] ,
         \s_mux2_signals[0][1][20] , \s_mux2_signals[0][1][19] ,
         \s_mux2_signals[0][1][18] , \s_mux2_signals[0][1][17] ,
         \s_mux2_signals[0][1][16] , \s_mux2_signals[0][1][15] ,
         \s_mux2_signals[0][1][14] , \s_mux2_signals[0][1][13] ,
         \s_mux2_signals[0][1][12] , \s_mux2_signals[0][1][11] ,
         \s_mux2_signals[0][1][10] , \s_mux2_signals[0][1][9] ,
         \s_mux2_signals[0][1][8] , \s_mux2_signals[0][1][7] ,
         \s_mux2_signals[0][1][6] , \s_mux2_signals[0][1][5] ,
         \s_mux2_signals[0][1][4] , \s_mux2_signals[0][1][3] ,
         \s_mux2_signals[0][1][2] , \s_mux2_signals[0][1][1] ,
         \s_mux2_signals[0][1][0] , \s_mux2_signals[0][2][31] ,
         \s_mux2_signals[0][2][30] , \s_mux2_signals[0][2][29] ,
         \s_mux2_signals[0][2][28] , \s_mux2_signals[0][2][27] ,
         \s_mux2_signals[0][2][26] , \s_mux2_signals[0][2][25] ,
         \s_mux2_signals[0][2][24] , \s_mux2_signals[0][2][23] ,
         \s_mux2_signals[0][2][22] , \s_mux2_signals[0][2][21] ,
         \s_mux2_signals[0][2][20] , \s_mux2_signals[0][2][19] ,
         \s_mux2_signals[0][2][18] , \s_mux2_signals[0][2][17] ,
         \s_mux2_signals[0][2][16] , \s_mux2_signals[0][2][15] ,
         \s_mux2_signals[0][2][14] , \s_mux2_signals[0][2][13] ,
         \s_mux2_signals[0][2][12] , \s_mux2_signals[0][2][11] ,
         \s_mux2_signals[0][2][10] , \s_mux2_signals[0][2][9] ,
         \s_mux2_signals[0][2][8] , \s_mux2_signals[0][2][7] ,
         \s_mux2_signals[0][2][6] , \s_mux2_signals[0][2][5] ,
         \s_mux2_signals[0][2][4] , \s_mux2_signals[0][2][3] ,
         \s_mux2_signals[0][2][2] , \s_mux2_signals[0][2][1] ,
         \s_mux2_signals[0][2][0] , \s_mux2_signals[0][3][31] ,
         \s_mux2_signals[0][3][30] , \s_mux2_signals[0][3][29] ,
         \s_mux2_signals[0][3][28] , \s_mux2_signals[0][3][27] ,
         \s_mux2_signals[0][3][26] , \s_mux2_signals[0][3][25] ,
         \s_mux2_signals[0][3][24] , \s_mux2_signals[0][3][23] ,
         \s_mux2_signals[0][3][22] , \s_mux2_signals[0][3][21] ,
         \s_mux2_signals[0][3][20] , \s_mux2_signals[0][3][19] ,
         \s_mux2_signals[0][3][18] , \s_mux2_signals[0][3][17] ,
         \s_mux2_signals[0][3][16] , \s_mux2_signals[0][3][15] ,
         \s_mux2_signals[0][3][14] , \s_mux2_signals[0][3][13] ,
         \s_mux2_signals[0][3][12] , \s_mux2_signals[0][3][11] ,
         \s_mux2_signals[0][3][10] , \s_mux2_signals[0][3][9] ,
         \s_mux2_signals[0][3][8] , \s_mux2_signals[0][3][7] ,
         \s_mux2_signals[0][3][6] , \s_mux2_signals[0][3][5] ,
         \s_mux2_signals[0][3][4] , \s_mux2_signals[0][3][3] ,
         \s_mux2_signals[0][3][2] , \s_mux2_signals[0][3][1] ,
         \s_mux2_signals[0][3][0] , \s_mux2_signals[0][4][31] ,
         \s_mux2_signals[0][4][30] , \s_mux2_signals[0][4][29] ,
         \s_mux2_signals[0][4][28] , \s_mux2_signals[0][4][27] ,
         \s_mux2_signals[0][4][26] , \s_mux2_signals[0][4][25] ,
         \s_mux2_signals[0][4][24] , \s_mux2_signals[0][4][23] ,
         \s_mux2_signals[0][4][22] , \s_mux2_signals[0][4][21] ,
         \s_mux2_signals[0][4][20] , \s_mux2_signals[0][4][19] ,
         \s_mux2_signals[0][4][18] , \s_mux2_signals[0][4][17] ,
         \s_mux2_signals[0][4][16] , \s_mux2_signals[0][4][15] ,
         \s_mux2_signals[0][4][14] , \s_mux2_signals[0][4][13] ,
         \s_mux2_signals[0][4][12] , \s_mux2_signals[0][4][11] ,
         \s_mux2_signals[0][4][10] , \s_mux2_signals[0][4][9] ,
         \s_mux2_signals[0][4][8] , \s_mux2_signals[0][4][7] ,
         \s_mux2_signals[0][4][6] , \s_mux2_signals[0][4][5] ,
         \s_mux2_signals[0][4][4] , \s_mux2_signals[0][4][3] ,
         \s_mux2_signals[0][4][2] , \s_mux2_signals[0][4][1] ,
         \s_mux2_signals[0][4][0] , \s_mux2_signals[0][5][31] ,
         \s_mux2_signals[0][5][30] , \s_mux2_signals[0][5][29] ,
         \s_mux2_signals[0][5][28] , \s_mux2_signals[0][5][27] ,
         \s_mux2_signals[0][5][26] , \s_mux2_signals[0][5][25] ,
         \s_mux2_signals[0][5][24] , \s_mux2_signals[0][5][23] ,
         \s_mux2_signals[0][5][22] , \s_mux2_signals[0][5][21] ,
         \s_mux2_signals[0][5][20] , \s_mux2_signals[0][5][19] ,
         \s_mux2_signals[0][5][18] , \s_mux2_signals[0][5][17] ,
         \s_mux2_signals[0][5][16] , \s_mux2_signals[0][5][15] ,
         \s_mux2_signals[0][5][14] , \s_mux2_signals[0][5][13] ,
         \s_mux2_signals[0][5][12] , \s_mux2_signals[0][5][11] ,
         \s_mux2_signals[0][5][10] , \s_mux2_signals[0][5][9] ,
         \s_mux2_signals[0][5][8] , \s_mux2_signals[0][5][7] ,
         \s_mux2_signals[0][5][6] , \s_mux2_signals[0][5][5] ,
         \s_mux2_signals[0][5][4] , \s_mux2_signals[0][5][3] ,
         \s_mux2_signals[0][5][2] , \s_mux2_signals[0][5][1] ,
         \s_mux2_signals[0][5][0] , \s_mux2_signals[0][6][31] ,
         \s_mux2_signals[0][6][30] , \s_mux2_signals[0][6][29] ,
         \s_mux2_signals[0][6][28] , \s_mux2_signals[0][6][27] ,
         \s_mux2_signals[0][6][26] , \s_mux2_signals[0][6][25] ,
         \s_mux2_signals[0][6][24] , \s_mux2_signals[0][6][23] ,
         \s_mux2_signals[0][6][22] , \s_mux2_signals[0][6][21] ,
         \s_mux2_signals[0][6][20] , \s_mux2_signals[0][6][19] ,
         \s_mux2_signals[0][6][18] , \s_mux2_signals[0][6][17] ,
         \s_mux2_signals[0][6][16] , \s_mux2_signals[0][6][15] ,
         \s_mux2_signals[0][6][14] , \s_mux2_signals[0][6][13] ,
         \s_mux2_signals[0][6][12] , \s_mux2_signals[0][6][11] ,
         \s_mux2_signals[0][6][10] , \s_mux2_signals[0][6][9] ,
         \s_mux2_signals[0][6][8] , \s_mux2_signals[0][6][7] ,
         \s_mux2_signals[0][6][6] , \s_mux2_signals[0][6][5] ,
         \s_mux2_signals[0][6][4] , \s_mux2_signals[0][6][3] ,
         \s_mux2_signals[0][6][2] , \s_mux2_signals[0][6][1] ,
         \s_mux2_signals[0][6][0] , \s_mux2_signals[0][7][31] ,
         \s_mux2_signals[0][7][30] , \s_mux2_signals[0][7][29] ,
         \s_mux2_signals[0][7][28] , \s_mux2_signals[0][7][27] ,
         \s_mux2_signals[0][7][26] , \s_mux2_signals[0][7][25] ,
         \s_mux2_signals[0][7][24] , \s_mux2_signals[0][7][23] ,
         \s_mux2_signals[0][7][22] , \s_mux2_signals[0][7][21] ,
         \s_mux2_signals[0][7][20] , \s_mux2_signals[0][7][19] ,
         \s_mux2_signals[0][7][18] , \s_mux2_signals[0][7][17] ,
         \s_mux2_signals[0][7][16] , \s_mux2_signals[0][7][15] ,
         \s_mux2_signals[0][7][14] , \s_mux2_signals[0][7][13] ,
         \s_mux2_signals[0][7][12] , \s_mux2_signals[0][7][11] ,
         \s_mux2_signals[0][7][10] , \s_mux2_signals[0][7][9] ,
         \s_mux2_signals[0][7][8] , \s_mux2_signals[0][7][7] ,
         \s_mux2_signals[0][7][6] , \s_mux2_signals[0][7][5] ,
         \s_mux2_signals[0][7][4] , \s_mux2_signals[0][7][3] ,
         \s_mux2_signals[0][7][2] , \s_mux2_signals[0][7][1] ,
         \s_mux2_signals[0][7][0] , \s_mux2_signals[0][8][31] ,
         \s_mux2_signals[0][8][30] , \s_mux2_signals[0][8][29] ,
         \s_mux2_signals[0][8][28] , \s_mux2_signals[0][8][27] ,
         \s_mux2_signals[0][8][26] , \s_mux2_signals[0][8][25] ,
         \s_mux2_signals[0][8][24] , \s_mux2_signals[0][8][23] ,
         \s_mux2_signals[0][8][22] , \s_mux2_signals[0][8][21] ,
         \s_mux2_signals[0][8][20] , \s_mux2_signals[0][8][19] ,
         \s_mux2_signals[0][8][18] , \s_mux2_signals[0][8][17] ,
         \s_mux2_signals[0][8][16] , \s_mux2_signals[0][8][15] ,
         \s_mux2_signals[0][8][14] , \s_mux2_signals[0][8][13] ,
         \s_mux2_signals[0][8][12] , \s_mux2_signals[0][8][11] ,
         \s_mux2_signals[0][8][10] , \s_mux2_signals[0][8][9] ,
         \s_mux2_signals[0][8][8] , \s_mux2_signals[0][8][7] ,
         \s_mux2_signals[0][8][6] , \s_mux2_signals[0][8][5] ,
         \s_mux2_signals[0][8][4] , \s_mux2_signals[0][8][3] ,
         \s_mux2_signals[0][8][2] , \s_mux2_signals[0][8][1] ,
         \s_mux2_signals[0][8][0] , \s_mux2_signals[0][9][31] ,
         \s_mux2_signals[0][9][30] , \s_mux2_signals[0][9][29] ,
         \s_mux2_signals[0][9][28] , \s_mux2_signals[0][9][27] ,
         \s_mux2_signals[0][9][26] , \s_mux2_signals[0][9][25] ,
         \s_mux2_signals[0][9][24] , \s_mux2_signals[0][9][23] ,
         \s_mux2_signals[0][9][22] , \s_mux2_signals[0][9][21] ,
         \s_mux2_signals[0][9][20] , \s_mux2_signals[0][9][19] ,
         \s_mux2_signals[0][9][18] , \s_mux2_signals[0][9][17] ,
         \s_mux2_signals[0][9][16] , \s_mux2_signals[0][9][15] ,
         \s_mux2_signals[0][9][14] , \s_mux2_signals[0][9][13] ,
         \s_mux2_signals[0][9][12] , \s_mux2_signals[0][9][11] ,
         \s_mux2_signals[0][9][10] , \s_mux2_signals[0][9][9] ,
         \s_mux2_signals[0][9][8] , \s_mux2_signals[0][9][7] ,
         \s_mux2_signals[0][9][6] , \s_mux2_signals[0][9][5] ,
         \s_mux2_signals[0][9][4] , \s_mux2_signals[0][9][3] ,
         \s_mux2_signals[0][9][2] , \s_mux2_signals[0][9][1] ,
         \s_mux2_signals[0][9][0] , \s_mux2_signals[0][10][31] ,
         \s_mux2_signals[0][10][30] , \s_mux2_signals[0][10][29] ,
         \s_mux2_signals[0][10][28] , \s_mux2_signals[0][10][27] ,
         \s_mux2_signals[0][10][26] , \s_mux2_signals[0][10][25] ,
         \s_mux2_signals[0][10][24] , \s_mux2_signals[0][10][23] ,
         \s_mux2_signals[0][10][22] , \s_mux2_signals[0][10][21] ,
         \s_mux2_signals[0][10][20] , \s_mux2_signals[0][10][19] ,
         \s_mux2_signals[0][10][18] , \s_mux2_signals[0][10][17] ,
         \s_mux2_signals[0][10][16] , \s_mux2_signals[0][10][15] ,
         \s_mux2_signals[0][10][14] , \s_mux2_signals[0][10][13] ,
         \s_mux2_signals[0][10][12] , \s_mux2_signals[0][10][11] ,
         \s_mux2_signals[0][10][10] , \s_mux2_signals[0][10][9] ,
         \s_mux2_signals[0][10][8] , \s_mux2_signals[0][10][7] ,
         \s_mux2_signals[0][10][6] , \s_mux2_signals[0][10][5] ,
         \s_mux2_signals[0][10][4] , \s_mux2_signals[0][10][3] ,
         \s_mux2_signals[0][10][2] , \s_mux2_signals[0][10][1] ,
         \s_mux2_signals[0][10][0] , \s_mux2_signals[0][11][31] ,
         \s_mux2_signals[0][11][30] , \s_mux2_signals[0][11][29] ,
         \s_mux2_signals[0][11][28] , \s_mux2_signals[0][11][27] ,
         \s_mux2_signals[0][11][26] , \s_mux2_signals[0][11][25] ,
         \s_mux2_signals[0][11][24] , \s_mux2_signals[0][11][23] ,
         \s_mux2_signals[0][11][22] , \s_mux2_signals[0][11][21] ,
         \s_mux2_signals[0][11][20] , \s_mux2_signals[0][11][19] ,
         \s_mux2_signals[0][11][18] , \s_mux2_signals[0][11][17] ,
         \s_mux2_signals[0][11][16] , \s_mux2_signals[0][11][15] ,
         \s_mux2_signals[0][11][14] , \s_mux2_signals[0][11][13] ,
         \s_mux2_signals[0][11][12] , \s_mux2_signals[0][11][11] ,
         \s_mux2_signals[0][11][10] , \s_mux2_signals[0][11][9] ,
         \s_mux2_signals[0][11][8] , \s_mux2_signals[0][11][7] ,
         \s_mux2_signals[0][11][6] , \s_mux2_signals[0][11][5] ,
         \s_mux2_signals[0][11][4] , \s_mux2_signals[0][11][3] ,
         \s_mux2_signals[0][11][2] , \s_mux2_signals[0][11][1] ,
         \s_mux2_signals[0][11][0] , \s_mux2_signals[0][12][31] ,
         \s_mux2_signals[0][12][30] , \s_mux2_signals[0][12][29] ,
         \s_mux2_signals[0][12][28] , \s_mux2_signals[0][12][27] ,
         \s_mux2_signals[0][12][26] , \s_mux2_signals[0][12][25] ,
         \s_mux2_signals[0][12][24] , \s_mux2_signals[0][12][23] ,
         \s_mux2_signals[0][12][22] , \s_mux2_signals[0][12][21] ,
         \s_mux2_signals[0][12][20] , \s_mux2_signals[0][12][19] ,
         \s_mux2_signals[0][12][18] , \s_mux2_signals[0][12][17] ,
         \s_mux2_signals[0][12][16] , \s_mux2_signals[0][12][15] ,
         \s_mux2_signals[0][12][14] , \s_mux2_signals[0][12][13] ,
         \s_mux2_signals[0][12][12] , \s_mux2_signals[0][12][11] ,
         \s_mux2_signals[0][12][10] , \s_mux2_signals[0][12][9] ,
         \s_mux2_signals[0][12][8] , \s_mux2_signals[0][12][7] ,
         \s_mux2_signals[0][12][6] , \s_mux2_signals[0][12][5] ,
         \s_mux2_signals[0][12][4] , \s_mux2_signals[0][12][3] ,
         \s_mux2_signals[0][12][2] , \s_mux2_signals[0][12][1] ,
         \s_mux2_signals[0][12][0] , \s_mux2_signals[0][13][31] ,
         \s_mux2_signals[0][13][30] , \s_mux2_signals[0][13][29] ,
         \s_mux2_signals[0][13][28] , \s_mux2_signals[0][13][27] ,
         \s_mux2_signals[0][13][26] , \s_mux2_signals[0][13][25] ,
         \s_mux2_signals[0][13][24] , \s_mux2_signals[0][13][23] ,
         \s_mux2_signals[0][13][22] , \s_mux2_signals[0][13][21] ,
         \s_mux2_signals[0][13][20] , \s_mux2_signals[0][13][19] ,
         \s_mux2_signals[0][13][18] , \s_mux2_signals[0][13][17] ,
         \s_mux2_signals[0][13][16] , \s_mux2_signals[0][13][15] ,
         \s_mux2_signals[0][13][14] , \s_mux2_signals[0][13][13] ,
         \s_mux2_signals[0][13][12] , \s_mux2_signals[0][13][11] ,
         \s_mux2_signals[0][13][10] , \s_mux2_signals[0][13][9] ,
         \s_mux2_signals[0][13][8] , \s_mux2_signals[0][13][7] ,
         \s_mux2_signals[0][13][6] , \s_mux2_signals[0][13][5] ,
         \s_mux2_signals[0][13][4] , \s_mux2_signals[0][13][3] ,
         \s_mux2_signals[0][13][2] , \s_mux2_signals[0][13][1] ,
         \s_mux2_signals[0][13][0] , \s_mux2_signals[0][14][31] ,
         \s_mux2_signals[0][14][30] , \s_mux2_signals[0][14][29] ,
         \s_mux2_signals[0][14][28] , \s_mux2_signals[0][14][27] ,
         \s_mux2_signals[0][14][26] , \s_mux2_signals[0][14][25] ,
         \s_mux2_signals[0][14][24] , \s_mux2_signals[0][14][23] ,
         \s_mux2_signals[0][14][22] , \s_mux2_signals[0][14][21] ,
         \s_mux2_signals[0][14][20] , \s_mux2_signals[0][14][19] ,
         \s_mux2_signals[0][14][18] , \s_mux2_signals[0][14][17] ,
         \s_mux2_signals[0][14][16] , \s_mux2_signals[0][14][15] ,
         \s_mux2_signals[0][14][14] , \s_mux2_signals[0][14][13] ,
         \s_mux2_signals[0][14][12] , \s_mux2_signals[0][14][11] ,
         \s_mux2_signals[0][14][10] , \s_mux2_signals[0][14][9] ,
         \s_mux2_signals[0][14][8] , \s_mux2_signals[0][14][7] ,
         \s_mux2_signals[0][14][6] , \s_mux2_signals[0][14][5] ,
         \s_mux2_signals[0][14][4] , \s_mux2_signals[0][14][3] ,
         \s_mux2_signals[0][14][2] , \s_mux2_signals[0][14][1] ,
         \s_mux2_signals[0][14][0] , \s_mux2_signals[0][15][31] ,
         \s_mux2_signals[0][15][30] , \s_mux2_signals[0][15][29] ,
         \s_mux2_signals[0][15][28] , \s_mux2_signals[0][15][27] ,
         \s_mux2_signals[0][15][26] , \s_mux2_signals[0][15][25] ,
         \s_mux2_signals[0][15][24] , \s_mux2_signals[0][15][23] ,
         \s_mux2_signals[0][15][22] , \s_mux2_signals[0][15][21] ,
         \s_mux2_signals[0][15][20] , \s_mux2_signals[0][15][19] ,
         \s_mux2_signals[0][15][18] , \s_mux2_signals[0][15][17] ,
         \s_mux2_signals[0][15][16] , \s_mux2_signals[0][15][15] ,
         \s_mux2_signals[0][15][14] , \s_mux2_signals[0][15][13] ,
         \s_mux2_signals[0][15][12] , \s_mux2_signals[0][15][11] ,
         \s_mux2_signals[0][15][10] , \s_mux2_signals[0][15][9] ,
         \s_mux2_signals[0][15][8] , \s_mux2_signals[0][15][7] ,
         \s_mux2_signals[0][15][6] , \s_mux2_signals[0][15][5] ,
         \s_mux2_signals[0][15][4] , \s_mux2_signals[0][15][3] ,
         \s_mux2_signals[0][15][2] , \s_mux2_signals[0][15][1] ,
         \s_mux2_signals[0][15][0] , \s_mux2_signals[0][16][31] ,
         \s_mux2_signals[0][16][30] , \s_mux2_signals[0][16][29] ,
         \s_mux2_signals[0][16][28] , \s_mux2_signals[0][16][27] ,
         \s_mux2_signals[0][16][26] , \s_mux2_signals[0][16][25] ,
         \s_mux2_signals[0][16][24] , \s_mux2_signals[0][16][23] ,
         \s_mux2_signals[0][16][22] , \s_mux2_signals[0][16][21] ,
         \s_mux2_signals[0][16][20] , \s_mux2_signals[0][16][19] ,
         \s_mux2_signals[0][16][18] , \s_mux2_signals[0][16][17] ,
         \s_mux2_signals[0][16][16] , \s_mux2_signals[0][16][15] ,
         \s_mux2_signals[0][16][14] , \s_mux2_signals[0][16][13] ,
         \s_mux2_signals[0][16][12] , \s_mux2_signals[0][16][11] ,
         \s_mux2_signals[0][16][10] , \s_mux2_signals[0][16][9] ,
         \s_mux2_signals[0][16][8] , \s_mux2_signals[0][16][7] ,
         \s_mux2_signals[0][16][6] , \s_mux2_signals[0][16][5] ,
         \s_mux2_signals[0][16][4] , \s_mux2_signals[0][16][3] ,
         \s_mux2_signals[0][16][2] , \s_mux2_signals[0][16][1] ,
         \s_mux2_signals[0][16][0] , \s_mux2_signals[0][17][31] ,
         \s_mux2_signals[0][17][30] , \s_mux2_signals[0][17][29] ,
         \s_mux2_signals[0][17][28] , \s_mux2_signals[0][17][27] ,
         \s_mux2_signals[0][17][26] , \s_mux2_signals[0][17][25] ,
         \s_mux2_signals[0][17][24] , \s_mux2_signals[0][17][23] ,
         \s_mux2_signals[0][17][22] , \s_mux2_signals[0][17][21] ,
         \s_mux2_signals[0][17][20] , \s_mux2_signals[0][17][19] ,
         \s_mux2_signals[0][17][18] , \s_mux2_signals[0][17][17] ,
         \s_mux2_signals[0][17][16] , \s_mux2_signals[0][17][15] ,
         \s_mux2_signals[0][17][14] , \s_mux2_signals[0][17][13] ,
         \s_mux2_signals[0][17][12] , \s_mux2_signals[0][17][11] ,
         \s_mux2_signals[0][17][10] , \s_mux2_signals[0][17][9] ,
         \s_mux2_signals[0][17][8] , \s_mux2_signals[0][17][7] ,
         \s_mux2_signals[0][17][6] , \s_mux2_signals[0][17][5] ,
         \s_mux2_signals[0][17][4] , \s_mux2_signals[0][17][3] ,
         \s_mux2_signals[0][17][2] , \s_mux2_signals[0][17][1] ,
         \s_mux2_signals[0][17][0] , \s_mux2_signals[0][18][31] ,
         \s_mux2_signals[0][18][30] , \s_mux2_signals[0][18][29] ,
         \s_mux2_signals[0][18][28] , \s_mux2_signals[0][18][27] ,
         \s_mux2_signals[0][18][26] , \s_mux2_signals[0][18][25] ,
         \s_mux2_signals[0][18][24] , \s_mux2_signals[0][18][23] ,
         \s_mux2_signals[0][18][22] , \s_mux2_signals[0][18][21] ,
         \s_mux2_signals[0][18][20] , \s_mux2_signals[0][18][19] ,
         \s_mux2_signals[0][18][18] , \s_mux2_signals[0][18][17] ,
         \s_mux2_signals[0][18][16] , \s_mux2_signals[0][18][15] ,
         \s_mux2_signals[0][18][14] , \s_mux2_signals[0][18][13] ,
         \s_mux2_signals[0][18][12] , \s_mux2_signals[0][18][11] ,
         \s_mux2_signals[0][18][10] , \s_mux2_signals[0][18][9] ,
         \s_mux2_signals[0][18][8] , \s_mux2_signals[0][18][7] ,
         \s_mux2_signals[0][18][6] , \s_mux2_signals[0][18][5] ,
         \s_mux2_signals[0][18][4] , \s_mux2_signals[0][18][3] ,
         \s_mux2_signals[0][18][2] , \s_mux2_signals[0][18][1] ,
         \s_mux2_signals[0][18][0] , \s_mux2_signals[0][19][31] ,
         \s_mux2_signals[0][19][30] , \s_mux2_signals[0][19][29] ,
         \s_mux2_signals[0][19][28] , \s_mux2_signals[0][19][27] ,
         \s_mux2_signals[0][19][26] , \s_mux2_signals[0][19][25] ,
         \s_mux2_signals[0][19][24] , \s_mux2_signals[0][19][23] ,
         \s_mux2_signals[0][19][22] , \s_mux2_signals[0][19][21] ,
         \s_mux2_signals[0][19][20] , \s_mux2_signals[0][19][19] ,
         \s_mux2_signals[0][19][18] , \s_mux2_signals[0][19][17] ,
         \s_mux2_signals[0][19][16] , \s_mux2_signals[0][19][15] ,
         \s_mux2_signals[0][19][14] , \s_mux2_signals[0][19][13] ,
         \s_mux2_signals[0][19][12] , \s_mux2_signals[0][19][11] ,
         \s_mux2_signals[0][19][10] , \s_mux2_signals[0][19][9] ,
         \s_mux2_signals[0][19][8] , \s_mux2_signals[0][19][7] ,
         \s_mux2_signals[0][19][6] , \s_mux2_signals[0][19][5] ,
         \s_mux2_signals[0][19][4] , \s_mux2_signals[0][19][3] ,
         \s_mux2_signals[0][19][2] , \s_mux2_signals[0][19][1] ,
         \s_mux2_signals[0][19][0] , \s_mux2_signals[0][20][31] ,
         \s_mux2_signals[0][20][30] , \s_mux2_signals[0][20][29] ,
         \s_mux2_signals[0][20][28] , \s_mux2_signals[0][20][27] ,
         \s_mux2_signals[0][20][26] , \s_mux2_signals[0][20][25] ,
         \s_mux2_signals[0][20][24] , \s_mux2_signals[0][20][23] ,
         \s_mux2_signals[0][20][22] , \s_mux2_signals[0][20][21] ,
         \s_mux2_signals[0][20][20] , \s_mux2_signals[0][20][19] ,
         \s_mux2_signals[0][20][18] , \s_mux2_signals[0][20][17] ,
         \s_mux2_signals[0][20][16] , \s_mux2_signals[0][20][15] ,
         \s_mux2_signals[0][20][14] , \s_mux2_signals[0][20][13] ,
         \s_mux2_signals[0][20][12] , \s_mux2_signals[0][20][11] ,
         \s_mux2_signals[0][20][10] , \s_mux2_signals[0][20][9] ,
         \s_mux2_signals[0][20][8] , \s_mux2_signals[0][20][7] ,
         \s_mux2_signals[0][20][6] , \s_mux2_signals[0][20][5] ,
         \s_mux2_signals[0][20][4] , \s_mux2_signals[0][20][3] ,
         \s_mux2_signals[0][20][2] , \s_mux2_signals[0][20][1] ,
         \s_mux2_signals[0][20][0] , \s_mux2_signals[0][21][31] ,
         \s_mux2_signals[0][21][30] , \s_mux2_signals[0][21][29] ,
         \s_mux2_signals[0][21][28] , \s_mux2_signals[0][21][27] ,
         \s_mux2_signals[0][21][26] , \s_mux2_signals[0][21][25] ,
         \s_mux2_signals[0][21][24] , \s_mux2_signals[0][21][23] ,
         \s_mux2_signals[0][21][22] , \s_mux2_signals[0][21][21] ,
         \s_mux2_signals[0][21][20] , \s_mux2_signals[0][21][19] ,
         \s_mux2_signals[0][21][18] , \s_mux2_signals[0][21][17] ,
         \s_mux2_signals[0][21][16] , \s_mux2_signals[0][21][15] ,
         \s_mux2_signals[0][21][14] , \s_mux2_signals[0][21][13] ,
         \s_mux2_signals[0][21][12] , \s_mux2_signals[0][21][11] ,
         \s_mux2_signals[0][21][10] , \s_mux2_signals[0][21][9] ,
         \s_mux2_signals[0][21][8] , \s_mux2_signals[0][21][7] ,
         \s_mux2_signals[0][21][6] , \s_mux2_signals[0][21][5] ,
         \s_mux2_signals[0][21][4] , \s_mux2_signals[0][21][3] ,
         \s_mux2_signals[0][21][2] , \s_mux2_signals[0][21][1] ,
         \s_mux2_signals[0][21][0] , \s_mux2_signals[0][22][31] ,
         \s_mux2_signals[0][22][30] , \s_mux2_signals[0][22][29] ,
         \s_mux2_signals[0][22][28] , \s_mux2_signals[0][22][27] ,
         \s_mux2_signals[0][22][26] , \s_mux2_signals[0][22][25] ,
         \s_mux2_signals[0][22][24] , \s_mux2_signals[0][22][23] ,
         \s_mux2_signals[0][22][22] , \s_mux2_signals[0][22][21] ,
         \s_mux2_signals[0][22][20] , \s_mux2_signals[0][22][19] ,
         \s_mux2_signals[0][22][18] , \s_mux2_signals[0][22][17] ,
         \s_mux2_signals[0][22][16] , \s_mux2_signals[0][22][15] ,
         \s_mux2_signals[0][22][14] , \s_mux2_signals[0][22][13] ,
         \s_mux2_signals[0][22][12] , \s_mux2_signals[0][22][11] ,
         \s_mux2_signals[0][22][10] , \s_mux2_signals[0][22][9] ,
         \s_mux2_signals[0][22][8] , \s_mux2_signals[0][22][7] ,
         \s_mux2_signals[0][22][6] , \s_mux2_signals[0][22][5] ,
         \s_mux2_signals[0][22][4] , \s_mux2_signals[0][22][3] ,
         \s_mux2_signals[0][22][2] , \s_mux2_signals[0][22][1] ,
         \s_mux2_signals[0][22][0] , \s_mux2_signals[0][23][31] ,
         \s_mux2_signals[0][23][30] , \s_mux2_signals[0][23][29] ,
         \s_mux2_signals[0][23][28] , \s_mux2_signals[0][23][27] ,
         \s_mux2_signals[0][23][26] , \s_mux2_signals[0][23][25] ,
         \s_mux2_signals[0][23][24] , \s_mux2_signals[0][23][23] ,
         \s_mux2_signals[0][23][22] , \s_mux2_signals[0][23][21] ,
         \s_mux2_signals[0][23][20] , \s_mux2_signals[0][23][19] ,
         \s_mux2_signals[0][23][18] , \s_mux2_signals[0][23][17] ,
         \s_mux2_signals[0][23][16] , \s_mux2_signals[0][23][15] ,
         \s_mux2_signals[0][23][14] , \s_mux2_signals[0][23][13] ,
         \s_mux2_signals[0][23][12] , \s_mux2_signals[0][23][11] ,
         \s_mux2_signals[0][23][10] , \s_mux2_signals[0][23][9] ,
         \s_mux2_signals[0][23][8] , \s_mux2_signals[0][23][7] ,
         \s_mux2_signals[0][23][6] , \s_mux2_signals[0][23][5] ,
         \s_mux2_signals[0][23][4] , \s_mux2_signals[0][23][3] ,
         \s_mux2_signals[0][23][2] , \s_mux2_signals[0][23][1] ,
         \s_mux2_signals[0][23][0] , \s_mux2_signals[0][24][31] ,
         \s_mux2_signals[0][24][30] , \s_mux2_signals[0][24][29] ,
         \s_mux2_signals[0][24][28] , \s_mux2_signals[0][24][27] ,
         \s_mux2_signals[0][24][26] , \s_mux2_signals[0][24][25] ,
         \s_mux2_signals[0][24][24] , \s_mux2_signals[0][24][23] ,
         \s_mux2_signals[0][24][22] , \s_mux2_signals[0][24][21] ,
         \s_mux2_signals[0][24][20] , \s_mux2_signals[0][24][19] ,
         \s_mux2_signals[0][24][18] , \s_mux2_signals[0][24][17] ,
         \s_mux2_signals[0][24][16] , \s_mux2_signals[0][24][15] ,
         \s_mux2_signals[0][24][14] , \s_mux2_signals[0][24][13] ,
         \s_mux2_signals[0][24][12] , \s_mux2_signals[0][24][11] ,
         \s_mux2_signals[0][24][10] , \s_mux2_signals[0][24][9] ,
         \s_mux2_signals[0][24][8] , \s_mux2_signals[0][24][7] ,
         \s_mux2_signals[0][24][6] , \s_mux2_signals[0][24][5] ,
         \s_mux2_signals[0][24][4] , \s_mux2_signals[0][24][3] ,
         \s_mux2_signals[0][24][2] , \s_mux2_signals[0][24][1] ,
         \s_mux2_signals[0][24][0] , \s_mux2_signals[0][25][31] ,
         \s_mux2_signals[0][25][30] , \s_mux2_signals[0][25][29] ,
         \s_mux2_signals[0][25][28] , \s_mux2_signals[0][25][27] ,
         \s_mux2_signals[0][25][26] , \s_mux2_signals[0][25][25] ,
         \s_mux2_signals[0][25][24] , \s_mux2_signals[0][25][23] ,
         \s_mux2_signals[0][25][22] , \s_mux2_signals[0][25][21] ,
         \s_mux2_signals[0][25][20] , \s_mux2_signals[0][25][19] ,
         \s_mux2_signals[0][25][18] , \s_mux2_signals[0][25][17] ,
         \s_mux2_signals[0][25][16] , \s_mux2_signals[0][25][15] ,
         \s_mux2_signals[0][25][14] , \s_mux2_signals[0][25][13] ,
         \s_mux2_signals[0][25][12] , \s_mux2_signals[0][25][11] ,
         \s_mux2_signals[0][25][10] , \s_mux2_signals[0][25][9] ,
         \s_mux2_signals[0][25][8] , \s_mux2_signals[0][25][7] ,
         \s_mux2_signals[0][25][6] , \s_mux2_signals[0][25][5] ,
         \s_mux2_signals[0][25][4] , \s_mux2_signals[0][25][3] ,
         \s_mux2_signals[0][25][2] , \s_mux2_signals[0][25][1] ,
         \s_mux2_signals[0][25][0] , \s_mux2_signals[0][26][31] ,
         \s_mux2_signals[0][26][30] , \s_mux2_signals[0][26][29] ,
         \s_mux2_signals[0][26][28] , \s_mux2_signals[0][26][27] ,
         \s_mux2_signals[0][26][26] , \s_mux2_signals[0][26][25] ,
         \s_mux2_signals[0][26][24] , \s_mux2_signals[0][26][23] ,
         \s_mux2_signals[0][26][22] , \s_mux2_signals[0][26][21] ,
         \s_mux2_signals[0][26][20] , \s_mux2_signals[0][26][19] ,
         \s_mux2_signals[0][26][18] , \s_mux2_signals[0][26][17] ,
         \s_mux2_signals[0][26][16] , \s_mux2_signals[0][26][15] ,
         \s_mux2_signals[0][26][14] , \s_mux2_signals[0][26][13] ,
         \s_mux2_signals[0][26][12] , \s_mux2_signals[0][26][11] ,
         \s_mux2_signals[0][26][10] , \s_mux2_signals[0][26][9] ,
         \s_mux2_signals[0][26][8] , \s_mux2_signals[0][26][7] ,
         \s_mux2_signals[0][26][6] , \s_mux2_signals[0][26][5] ,
         \s_mux2_signals[0][26][4] , \s_mux2_signals[0][26][3] ,
         \s_mux2_signals[0][26][2] , \s_mux2_signals[0][26][1] ,
         \s_mux2_signals[0][26][0] , \s_mux2_signals[0][27][31] ,
         \s_mux2_signals[0][27][30] , \s_mux2_signals[0][27][29] ,
         \s_mux2_signals[0][27][28] , \s_mux2_signals[0][27][27] ,
         \s_mux2_signals[0][27][26] , \s_mux2_signals[0][27][25] ,
         \s_mux2_signals[0][27][24] , \s_mux2_signals[0][27][23] ,
         \s_mux2_signals[0][27][22] , \s_mux2_signals[0][27][21] ,
         \s_mux2_signals[0][27][20] , \s_mux2_signals[0][27][19] ,
         \s_mux2_signals[0][27][18] , \s_mux2_signals[0][27][17] ,
         \s_mux2_signals[0][27][16] , \s_mux2_signals[0][27][15] ,
         \s_mux2_signals[0][27][14] , \s_mux2_signals[0][27][13] ,
         \s_mux2_signals[0][27][12] , \s_mux2_signals[0][27][11] ,
         \s_mux2_signals[0][27][10] , \s_mux2_signals[0][27][9] ,
         \s_mux2_signals[0][27][8] , \s_mux2_signals[0][27][7] ,
         \s_mux2_signals[0][27][6] , \s_mux2_signals[0][27][5] ,
         \s_mux2_signals[0][27][4] , \s_mux2_signals[0][27][3] ,
         \s_mux2_signals[0][27][2] , \s_mux2_signals[0][27][1] ,
         \s_mux2_signals[0][27][0] , \s_mux2_signals[0][28][31] ,
         \s_mux2_signals[0][28][30] , \s_mux2_signals[0][28][29] ,
         \s_mux2_signals[0][28][28] , \s_mux2_signals[0][28][27] ,
         \s_mux2_signals[0][28][26] , \s_mux2_signals[0][28][25] ,
         \s_mux2_signals[0][28][24] , \s_mux2_signals[0][28][23] ,
         \s_mux2_signals[0][28][22] , \s_mux2_signals[0][28][21] ,
         \s_mux2_signals[0][28][20] , \s_mux2_signals[0][28][19] ,
         \s_mux2_signals[0][28][18] , \s_mux2_signals[0][28][17] ,
         \s_mux2_signals[0][28][16] , \s_mux2_signals[0][28][15] ,
         \s_mux2_signals[0][28][14] , \s_mux2_signals[0][28][13] ,
         \s_mux2_signals[0][28][12] , \s_mux2_signals[0][28][11] ,
         \s_mux2_signals[0][28][10] , \s_mux2_signals[0][28][9] ,
         \s_mux2_signals[0][28][8] , \s_mux2_signals[0][28][7] ,
         \s_mux2_signals[0][28][6] , \s_mux2_signals[0][28][5] ,
         \s_mux2_signals[0][28][4] , \s_mux2_signals[0][28][3] ,
         \s_mux2_signals[0][28][2] , \s_mux2_signals[0][28][1] ,
         \s_mux2_signals[0][28][0] , \s_mux2_signals[0][29][31] ,
         \s_mux2_signals[0][29][30] , \s_mux2_signals[0][29][29] ,
         \s_mux2_signals[0][29][28] , \s_mux2_signals[0][29][27] ,
         \s_mux2_signals[0][29][26] , \s_mux2_signals[0][29][25] ,
         \s_mux2_signals[0][29][24] , \s_mux2_signals[0][29][23] ,
         \s_mux2_signals[0][29][22] , \s_mux2_signals[0][29][21] ,
         \s_mux2_signals[0][29][20] , \s_mux2_signals[0][29][19] ,
         \s_mux2_signals[0][29][18] , \s_mux2_signals[0][29][17] ,
         \s_mux2_signals[0][29][16] , \s_mux2_signals[0][29][15] ,
         \s_mux2_signals[0][29][14] , \s_mux2_signals[0][29][13] ,
         \s_mux2_signals[0][29][12] , \s_mux2_signals[0][29][11] ,
         \s_mux2_signals[0][29][10] , \s_mux2_signals[0][29][9] ,
         \s_mux2_signals[0][29][8] , \s_mux2_signals[0][29][7] ,
         \s_mux2_signals[0][29][6] , \s_mux2_signals[0][29][5] ,
         \s_mux2_signals[0][29][4] , \s_mux2_signals[0][29][3] ,
         \s_mux2_signals[0][29][2] , \s_mux2_signals[0][29][1] ,
         \s_mux2_signals[0][29][0] , \s_mux2_signals[0][30][31] ,
         \s_mux2_signals[0][30][30] , \s_mux2_signals[0][30][29] ,
         \s_mux2_signals[0][30][28] , \s_mux2_signals[0][30][27] ,
         \s_mux2_signals[0][30][26] , \s_mux2_signals[0][30][25] ,
         \s_mux2_signals[0][30][24] , \s_mux2_signals[0][30][23] ,
         \s_mux2_signals[0][30][22] , \s_mux2_signals[0][30][21] ,
         \s_mux2_signals[0][30][20] , \s_mux2_signals[0][30][19] ,
         \s_mux2_signals[0][30][18] , \s_mux2_signals[0][30][17] ,
         \s_mux2_signals[0][30][16] , \s_mux2_signals[0][30][15] ,
         \s_mux2_signals[0][30][14] , \s_mux2_signals[0][30][13] ,
         \s_mux2_signals[0][30][12] , \s_mux2_signals[0][30][11] ,
         \s_mux2_signals[0][30][10] , \s_mux2_signals[0][30][9] ,
         \s_mux2_signals[0][30][8] , \s_mux2_signals[0][30][7] ,
         \s_mux2_signals[0][30][6] , \s_mux2_signals[0][30][5] ,
         \s_mux2_signals[0][30][4] , \s_mux2_signals[0][30][3] ,
         \s_mux2_signals[0][30][2] , \s_mux2_signals[0][30][1] ,
         \s_mux2_signals[0][30][0] , \s_mux2_signals[0][31][31] ,
         \s_mux2_signals[0][31][30] , \s_mux2_signals[0][31][29] ,
         \s_mux2_signals[0][31][28] , \s_mux2_signals[0][31][27] ,
         \s_mux2_signals[0][31][26] , \s_mux2_signals[0][31][25] ,
         \s_mux2_signals[0][31][24] , \s_mux2_signals[0][31][23] ,
         \s_mux2_signals[0][31][22] , \s_mux2_signals[0][31][21] ,
         \s_mux2_signals[0][31][20] , \s_mux2_signals[0][31][19] ,
         \s_mux2_signals[0][31][18] , \s_mux2_signals[0][31][17] ,
         \s_mux2_signals[0][31][16] , \s_mux2_signals[0][31][15] ,
         \s_mux2_signals[0][31][14] , \s_mux2_signals[0][31][13] ,
         \s_mux2_signals[0][31][12] , \s_mux2_signals[0][31][11] ,
         \s_mux2_signals[0][31][10] , \s_mux2_signals[0][31][9] ,
         \s_mux2_signals[0][31][8] , \s_mux2_signals[0][31][7] ,
         \s_mux2_signals[0][31][6] , \s_mux2_signals[0][31][5] ,
         \s_mux2_signals[0][31][4] , \s_mux2_signals[0][31][3] ,
         \s_mux2_signals[0][31][2] , \s_mux2_signals[0][31][1] ,
         \s_mux2_signals[0][31][0] , \s_mux2_signals[1][0][31] ,
         \s_mux2_signals[1][0][30] , \s_mux2_signals[1][0][29] ,
         \s_mux2_signals[1][0][28] , \s_mux2_signals[1][0][27] ,
         \s_mux2_signals[1][0][26] , \s_mux2_signals[1][0][25] ,
         \s_mux2_signals[1][0][24] , \s_mux2_signals[1][0][23] ,
         \s_mux2_signals[1][0][22] , \s_mux2_signals[1][0][21] ,
         \s_mux2_signals[1][0][20] , \s_mux2_signals[1][0][19] ,
         \s_mux2_signals[1][0][18] , \s_mux2_signals[1][0][17] ,
         \s_mux2_signals[1][0][16] , \s_mux2_signals[1][0][15] ,
         \s_mux2_signals[1][0][14] , \s_mux2_signals[1][0][13] ,
         \s_mux2_signals[1][0][12] , \s_mux2_signals[1][0][11] ,
         \s_mux2_signals[1][0][10] , \s_mux2_signals[1][0][9] ,
         \s_mux2_signals[1][0][8] , \s_mux2_signals[1][0][7] ,
         \s_mux2_signals[1][0][6] , \s_mux2_signals[1][0][5] ,
         \s_mux2_signals[1][0][4] , \s_mux2_signals[1][0][3] ,
         \s_mux2_signals[1][0][2] , \s_mux2_signals[1][0][1] ,
         \s_mux2_signals[1][0][0] , \s_mux2_signals[1][2][31] ,
         \s_mux2_signals[1][2][30] , \s_mux2_signals[1][2][29] ,
         \s_mux2_signals[1][2][28] , \s_mux2_signals[1][2][27] ,
         \s_mux2_signals[1][2][26] , \s_mux2_signals[1][2][25] ,
         \s_mux2_signals[1][2][24] , \s_mux2_signals[1][2][23] ,
         \s_mux2_signals[1][2][22] , \s_mux2_signals[1][2][21] ,
         \s_mux2_signals[1][2][20] , \s_mux2_signals[1][2][19] ,
         \s_mux2_signals[1][2][18] , \s_mux2_signals[1][2][17] ,
         \s_mux2_signals[1][2][16] , \s_mux2_signals[1][2][15] ,
         \s_mux2_signals[1][2][14] , \s_mux2_signals[1][2][13] ,
         \s_mux2_signals[1][2][12] , \s_mux2_signals[1][2][11] ,
         \s_mux2_signals[1][2][10] , \s_mux2_signals[1][2][9] ,
         \s_mux2_signals[1][2][8] , \s_mux2_signals[1][2][7] ,
         \s_mux2_signals[1][2][6] , \s_mux2_signals[1][2][5] ,
         \s_mux2_signals[1][2][4] , \s_mux2_signals[1][2][3] ,
         \s_mux2_signals[1][2][2] , \s_mux2_signals[1][2][1] ,
         \s_mux2_signals[1][2][0] , \s_mux2_signals[1][4][31] ,
         \s_mux2_signals[1][4][30] , \s_mux2_signals[1][4][29] ,
         \s_mux2_signals[1][4][28] , \s_mux2_signals[1][4][27] ,
         \s_mux2_signals[1][4][26] , \s_mux2_signals[1][4][25] ,
         \s_mux2_signals[1][4][24] , \s_mux2_signals[1][4][23] ,
         \s_mux2_signals[1][4][22] , \s_mux2_signals[1][4][21] ,
         \s_mux2_signals[1][4][20] , \s_mux2_signals[1][4][19] ,
         \s_mux2_signals[1][4][18] , \s_mux2_signals[1][4][17] ,
         \s_mux2_signals[1][4][16] , \s_mux2_signals[1][4][15] ,
         \s_mux2_signals[1][4][14] , \s_mux2_signals[1][4][13] ,
         \s_mux2_signals[1][4][12] , \s_mux2_signals[1][4][11] ,
         \s_mux2_signals[1][4][10] , \s_mux2_signals[1][4][9] ,
         \s_mux2_signals[1][4][8] , \s_mux2_signals[1][4][7] ,
         \s_mux2_signals[1][4][6] , \s_mux2_signals[1][4][5] ,
         \s_mux2_signals[1][4][4] , \s_mux2_signals[1][4][3] ,
         \s_mux2_signals[1][4][2] , \s_mux2_signals[1][4][1] ,
         \s_mux2_signals[1][4][0] , \s_mux2_signals[1][6][31] ,
         \s_mux2_signals[1][6][30] , \s_mux2_signals[1][6][29] ,
         \s_mux2_signals[1][6][28] , \s_mux2_signals[1][6][27] ,
         \s_mux2_signals[1][6][26] , \s_mux2_signals[1][6][25] ,
         \s_mux2_signals[1][6][24] , \s_mux2_signals[1][6][23] ,
         \s_mux2_signals[1][6][22] , \s_mux2_signals[1][6][21] ,
         \s_mux2_signals[1][6][20] , \s_mux2_signals[1][6][19] ,
         \s_mux2_signals[1][6][18] , \s_mux2_signals[1][6][17] ,
         \s_mux2_signals[1][6][16] , \s_mux2_signals[1][6][15] ,
         \s_mux2_signals[1][6][14] , \s_mux2_signals[1][6][13] ,
         \s_mux2_signals[1][6][12] , \s_mux2_signals[1][6][11] ,
         \s_mux2_signals[1][6][10] , \s_mux2_signals[1][6][9] ,
         \s_mux2_signals[1][6][8] , \s_mux2_signals[1][6][7] ,
         \s_mux2_signals[1][6][6] , \s_mux2_signals[1][6][5] ,
         \s_mux2_signals[1][6][4] , \s_mux2_signals[1][6][3] ,
         \s_mux2_signals[1][6][2] , \s_mux2_signals[1][6][1] ,
         \s_mux2_signals[1][6][0] , \s_mux2_signals[1][8][31] ,
         \s_mux2_signals[1][8][30] , \s_mux2_signals[1][8][29] ,
         \s_mux2_signals[1][8][28] , \s_mux2_signals[1][8][27] ,
         \s_mux2_signals[1][8][26] , \s_mux2_signals[1][8][25] ,
         \s_mux2_signals[1][8][24] , \s_mux2_signals[1][8][23] ,
         \s_mux2_signals[1][8][22] , \s_mux2_signals[1][8][21] ,
         \s_mux2_signals[1][8][20] , \s_mux2_signals[1][8][19] ,
         \s_mux2_signals[1][8][18] , \s_mux2_signals[1][8][17] ,
         \s_mux2_signals[1][8][16] , \s_mux2_signals[1][8][15] ,
         \s_mux2_signals[1][8][14] , \s_mux2_signals[1][8][13] ,
         \s_mux2_signals[1][8][12] , \s_mux2_signals[1][8][11] ,
         \s_mux2_signals[1][8][10] , \s_mux2_signals[1][8][9] ,
         \s_mux2_signals[1][8][8] , \s_mux2_signals[1][8][7] ,
         \s_mux2_signals[1][8][6] , \s_mux2_signals[1][8][5] ,
         \s_mux2_signals[1][8][4] , \s_mux2_signals[1][8][3] ,
         \s_mux2_signals[1][8][2] , \s_mux2_signals[1][8][1] ,
         \s_mux2_signals[1][8][0] , \s_mux2_signals[1][10][31] ,
         \s_mux2_signals[1][10][30] , \s_mux2_signals[1][10][29] ,
         \s_mux2_signals[1][10][28] , \s_mux2_signals[1][10][27] ,
         \s_mux2_signals[1][10][26] , \s_mux2_signals[1][10][25] ,
         \s_mux2_signals[1][10][24] , \s_mux2_signals[1][10][23] ,
         \s_mux2_signals[1][10][22] , \s_mux2_signals[1][10][21] ,
         \s_mux2_signals[1][10][20] , \s_mux2_signals[1][10][19] ,
         \s_mux2_signals[1][10][18] , \s_mux2_signals[1][10][17] ,
         \s_mux2_signals[1][10][16] , \s_mux2_signals[1][10][15] ,
         \s_mux2_signals[1][10][14] , \s_mux2_signals[1][10][13] ,
         \s_mux2_signals[1][10][12] , \s_mux2_signals[1][10][11] ,
         \s_mux2_signals[1][10][10] , \s_mux2_signals[1][10][9] ,
         \s_mux2_signals[1][10][8] , \s_mux2_signals[1][10][7] ,
         \s_mux2_signals[1][10][6] , \s_mux2_signals[1][10][5] ,
         \s_mux2_signals[1][10][4] , \s_mux2_signals[1][10][3] ,
         \s_mux2_signals[1][10][2] , \s_mux2_signals[1][10][1] ,
         \s_mux2_signals[1][10][0] , \s_mux2_signals[1][12][31] ,
         \s_mux2_signals[1][12][30] , \s_mux2_signals[1][12][29] ,
         \s_mux2_signals[1][12][28] , \s_mux2_signals[1][12][27] ,
         \s_mux2_signals[1][12][26] , \s_mux2_signals[1][12][25] ,
         \s_mux2_signals[1][12][24] , \s_mux2_signals[1][12][23] ,
         \s_mux2_signals[1][12][22] , \s_mux2_signals[1][12][21] ,
         \s_mux2_signals[1][12][20] , \s_mux2_signals[1][12][19] ,
         \s_mux2_signals[1][12][18] , \s_mux2_signals[1][12][17] ,
         \s_mux2_signals[1][12][16] , \s_mux2_signals[1][12][15] ,
         \s_mux2_signals[1][12][14] , \s_mux2_signals[1][12][13] ,
         \s_mux2_signals[1][12][12] , \s_mux2_signals[1][12][11] ,
         \s_mux2_signals[1][12][10] , \s_mux2_signals[1][12][9] ,
         \s_mux2_signals[1][12][8] , \s_mux2_signals[1][12][7] ,
         \s_mux2_signals[1][12][6] , \s_mux2_signals[1][12][5] ,
         \s_mux2_signals[1][12][4] , \s_mux2_signals[1][12][3] ,
         \s_mux2_signals[1][12][2] , \s_mux2_signals[1][12][1] ,
         \s_mux2_signals[1][12][0] , \s_mux2_signals[1][14][31] ,
         \s_mux2_signals[1][14][30] , \s_mux2_signals[1][14][29] ,
         \s_mux2_signals[1][14][28] , \s_mux2_signals[1][14][27] ,
         \s_mux2_signals[1][14][26] , \s_mux2_signals[1][14][25] ,
         \s_mux2_signals[1][14][24] , \s_mux2_signals[1][14][23] ,
         \s_mux2_signals[1][14][22] , \s_mux2_signals[1][14][21] ,
         \s_mux2_signals[1][14][20] , \s_mux2_signals[1][14][19] ,
         \s_mux2_signals[1][14][18] , \s_mux2_signals[1][14][17] ,
         \s_mux2_signals[1][14][16] , \s_mux2_signals[1][14][15] ,
         \s_mux2_signals[1][14][14] , \s_mux2_signals[1][14][13] ,
         \s_mux2_signals[1][14][12] , \s_mux2_signals[1][14][11] ,
         \s_mux2_signals[1][14][10] , \s_mux2_signals[1][14][9] ,
         \s_mux2_signals[1][14][8] , \s_mux2_signals[1][14][7] ,
         \s_mux2_signals[1][14][6] , \s_mux2_signals[1][14][5] ,
         \s_mux2_signals[1][14][4] , \s_mux2_signals[1][14][3] ,
         \s_mux2_signals[1][14][2] , \s_mux2_signals[1][14][1] ,
         \s_mux2_signals[1][14][0] , \s_mux2_signals[1][16][31] ,
         \s_mux2_signals[1][16][30] , \s_mux2_signals[1][16][29] ,
         \s_mux2_signals[1][16][28] , \s_mux2_signals[1][16][27] ,
         \s_mux2_signals[1][16][26] , \s_mux2_signals[1][16][25] ,
         \s_mux2_signals[1][16][24] , \s_mux2_signals[1][16][23] ,
         \s_mux2_signals[1][16][22] , \s_mux2_signals[1][16][21] ,
         \s_mux2_signals[1][16][20] , \s_mux2_signals[1][16][19] ,
         \s_mux2_signals[1][16][18] , \s_mux2_signals[1][16][17] ,
         \s_mux2_signals[1][16][16] , \s_mux2_signals[1][16][15] ,
         \s_mux2_signals[1][16][14] , \s_mux2_signals[1][16][13] ,
         \s_mux2_signals[1][16][12] , \s_mux2_signals[1][16][11] ,
         \s_mux2_signals[1][16][10] , \s_mux2_signals[1][16][9] ,
         \s_mux2_signals[1][16][8] , \s_mux2_signals[1][16][7] ,
         \s_mux2_signals[1][16][6] , \s_mux2_signals[1][16][5] ,
         \s_mux2_signals[1][16][4] , \s_mux2_signals[1][16][3] ,
         \s_mux2_signals[1][16][2] , \s_mux2_signals[1][16][1] ,
         \s_mux2_signals[1][16][0] , \s_mux2_signals[1][18][31] ,
         \s_mux2_signals[1][18][30] , \s_mux2_signals[1][18][29] ,
         \s_mux2_signals[1][18][28] , \s_mux2_signals[1][18][27] ,
         \s_mux2_signals[1][18][26] , \s_mux2_signals[1][18][25] ,
         \s_mux2_signals[1][18][24] , \s_mux2_signals[1][18][23] ,
         \s_mux2_signals[1][18][22] , \s_mux2_signals[1][18][21] ,
         \s_mux2_signals[1][18][20] , \s_mux2_signals[1][18][19] ,
         \s_mux2_signals[1][18][18] , \s_mux2_signals[1][18][17] ,
         \s_mux2_signals[1][18][16] , \s_mux2_signals[1][18][15] ,
         \s_mux2_signals[1][18][14] , \s_mux2_signals[1][18][13] ,
         \s_mux2_signals[1][18][12] , \s_mux2_signals[1][18][11] ,
         \s_mux2_signals[1][18][10] , \s_mux2_signals[1][18][9] ,
         \s_mux2_signals[1][18][8] , \s_mux2_signals[1][18][7] ,
         \s_mux2_signals[1][18][6] , \s_mux2_signals[1][18][5] ,
         \s_mux2_signals[1][18][4] , \s_mux2_signals[1][18][3] ,
         \s_mux2_signals[1][18][2] , \s_mux2_signals[1][18][1] ,
         \s_mux2_signals[1][18][0] , \s_mux2_signals[1][20][31] ,
         \s_mux2_signals[1][20][30] , \s_mux2_signals[1][20][29] ,
         \s_mux2_signals[1][20][28] , \s_mux2_signals[1][20][27] ,
         \s_mux2_signals[1][20][26] , \s_mux2_signals[1][20][25] ,
         \s_mux2_signals[1][20][24] , \s_mux2_signals[1][20][23] ,
         \s_mux2_signals[1][20][22] , \s_mux2_signals[1][20][21] ,
         \s_mux2_signals[1][20][20] , \s_mux2_signals[1][20][19] ,
         \s_mux2_signals[1][20][18] , \s_mux2_signals[1][20][17] ,
         \s_mux2_signals[1][20][16] , \s_mux2_signals[1][20][15] ,
         \s_mux2_signals[1][20][14] , \s_mux2_signals[1][20][13] ,
         \s_mux2_signals[1][20][12] , \s_mux2_signals[1][20][11] ,
         \s_mux2_signals[1][20][10] , \s_mux2_signals[1][20][9] ,
         \s_mux2_signals[1][20][8] , \s_mux2_signals[1][20][7] ,
         \s_mux2_signals[1][20][6] , \s_mux2_signals[1][20][5] ,
         \s_mux2_signals[1][20][4] , \s_mux2_signals[1][20][3] ,
         \s_mux2_signals[1][20][2] , \s_mux2_signals[1][20][1] ,
         \s_mux2_signals[1][20][0] , \s_mux2_signals[1][22][31] ,
         \s_mux2_signals[1][22][30] , \s_mux2_signals[1][22][29] ,
         \s_mux2_signals[1][22][28] , \s_mux2_signals[1][22][27] ,
         \s_mux2_signals[1][22][26] , \s_mux2_signals[1][22][25] ,
         \s_mux2_signals[1][22][24] , \s_mux2_signals[1][22][23] ,
         \s_mux2_signals[1][22][22] , \s_mux2_signals[1][22][21] ,
         \s_mux2_signals[1][22][20] , \s_mux2_signals[1][22][19] ,
         \s_mux2_signals[1][22][18] , \s_mux2_signals[1][22][17] ,
         \s_mux2_signals[1][22][16] , \s_mux2_signals[1][22][15] ,
         \s_mux2_signals[1][22][14] , \s_mux2_signals[1][22][13] ,
         \s_mux2_signals[1][22][12] , \s_mux2_signals[1][22][11] ,
         \s_mux2_signals[1][22][10] , \s_mux2_signals[1][22][9] ,
         \s_mux2_signals[1][22][8] , \s_mux2_signals[1][22][7] ,
         \s_mux2_signals[1][22][6] , \s_mux2_signals[1][22][5] ,
         \s_mux2_signals[1][22][4] , \s_mux2_signals[1][22][3] ,
         \s_mux2_signals[1][22][2] , \s_mux2_signals[1][22][1] ,
         \s_mux2_signals[1][22][0] , \s_mux2_signals[1][24][31] ,
         \s_mux2_signals[1][24][30] , \s_mux2_signals[1][24][29] ,
         \s_mux2_signals[1][24][28] , \s_mux2_signals[1][24][27] ,
         \s_mux2_signals[1][24][26] , \s_mux2_signals[1][24][25] ,
         \s_mux2_signals[1][24][24] , \s_mux2_signals[1][24][23] ,
         \s_mux2_signals[1][24][22] , \s_mux2_signals[1][24][21] ,
         \s_mux2_signals[1][24][20] , \s_mux2_signals[1][24][19] ,
         \s_mux2_signals[1][24][18] , \s_mux2_signals[1][24][17] ,
         \s_mux2_signals[1][24][16] , \s_mux2_signals[1][24][15] ,
         \s_mux2_signals[1][24][14] , \s_mux2_signals[1][24][13] ,
         \s_mux2_signals[1][24][12] , \s_mux2_signals[1][24][11] ,
         \s_mux2_signals[1][24][10] , \s_mux2_signals[1][24][9] ,
         \s_mux2_signals[1][24][8] , \s_mux2_signals[1][24][7] ,
         \s_mux2_signals[1][24][6] , \s_mux2_signals[1][24][5] ,
         \s_mux2_signals[1][24][4] , \s_mux2_signals[1][24][3] ,
         \s_mux2_signals[1][24][2] , \s_mux2_signals[1][24][1] ,
         \s_mux2_signals[1][24][0] , \s_mux2_signals[1][26][31] ,
         \s_mux2_signals[1][26][30] , \s_mux2_signals[1][26][29] ,
         \s_mux2_signals[1][26][28] , \s_mux2_signals[1][26][27] ,
         \s_mux2_signals[1][26][26] , \s_mux2_signals[1][26][25] ,
         \s_mux2_signals[1][26][24] , \s_mux2_signals[1][26][23] ,
         \s_mux2_signals[1][26][22] , \s_mux2_signals[1][26][21] ,
         \s_mux2_signals[1][26][20] , \s_mux2_signals[1][26][19] ,
         \s_mux2_signals[1][26][18] , \s_mux2_signals[1][26][17] ,
         \s_mux2_signals[1][26][16] , \s_mux2_signals[1][26][15] ,
         \s_mux2_signals[1][26][14] , \s_mux2_signals[1][26][13] ,
         \s_mux2_signals[1][26][12] , \s_mux2_signals[1][26][11] ,
         \s_mux2_signals[1][26][10] , \s_mux2_signals[1][26][9] ,
         \s_mux2_signals[1][26][8] , \s_mux2_signals[1][26][7] ,
         \s_mux2_signals[1][26][6] , \s_mux2_signals[1][26][5] ,
         \s_mux2_signals[1][26][4] , \s_mux2_signals[1][26][3] ,
         \s_mux2_signals[1][26][2] , \s_mux2_signals[1][26][1] ,
         \s_mux2_signals[1][26][0] , \s_mux2_signals[1][28][31] ,
         \s_mux2_signals[1][28][30] , \s_mux2_signals[1][28][29] ,
         \s_mux2_signals[1][28][28] , \s_mux2_signals[1][28][27] ,
         \s_mux2_signals[1][28][26] , \s_mux2_signals[1][28][25] ,
         \s_mux2_signals[1][28][24] , \s_mux2_signals[1][28][23] ,
         \s_mux2_signals[1][28][22] , \s_mux2_signals[1][28][21] ,
         \s_mux2_signals[1][28][20] , \s_mux2_signals[1][28][19] ,
         \s_mux2_signals[1][28][18] , \s_mux2_signals[1][28][17] ,
         \s_mux2_signals[1][28][16] , \s_mux2_signals[1][28][15] ,
         \s_mux2_signals[1][28][14] , \s_mux2_signals[1][28][13] ,
         \s_mux2_signals[1][28][12] , \s_mux2_signals[1][28][11] ,
         \s_mux2_signals[1][28][10] , \s_mux2_signals[1][28][9] ,
         \s_mux2_signals[1][28][8] , \s_mux2_signals[1][28][7] ,
         \s_mux2_signals[1][28][6] , \s_mux2_signals[1][28][5] ,
         \s_mux2_signals[1][28][4] , \s_mux2_signals[1][28][3] ,
         \s_mux2_signals[1][28][2] , \s_mux2_signals[1][28][1] ,
         \s_mux2_signals[1][28][0] , \s_mux2_signals[1][30][31] ,
         \s_mux2_signals[1][30][30] , \s_mux2_signals[1][30][29] ,
         \s_mux2_signals[1][30][28] , \s_mux2_signals[1][30][27] ,
         \s_mux2_signals[1][30][26] , \s_mux2_signals[1][30][25] ,
         \s_mux2_signals[1][30][24] , \s_mux2_signals[1][30][23] ,
         \s_mux2_signals[1][30][22] , \s_mux2_signals[1][30][21] ,
         \s_mux2_signals[1][30][20] , \s_mux2_signals[1][30][19] ,
         \s_mux2_signals[1][30][18] , \s_mux2_signals[1][30][17] ,
         \s_mux2_signals[1][30][16] , \s_mux2_signals[1][30][15] ,
         \s_mux2_signals[1][30][14] , \s_mux2_signals[1][30][13] ,
         \s_mux2_signals[1][30][12] , \s_mux2_signals[1][30][11] ,
         \s_mux2_signals[1][30][10] , \s_mux2_signals[1][30][9] ,
         \s_mux2_signals[1][30][8] , \s_mux2_signals[1][30][7] ,
         \s_mux2_signals[1][30][6] , \s_mux2_signals[1][30][5] ,
         \s_mux2_signals[1][30][4] , \s_mux2_signals[1][30][3] ,
         \s_mux2_signals[1][30][2] , \s_mux2_signals[1][30][1] ,
         \s_mux2_signals[1][30][0] , \s_mux2_signals[2][0][31] ,
         \s_mux2_signals[2][0][30] , \s_mux2_signals[2][0][29] ,
         \s_mux2_signals[2][0][28] , \s_mux2_signals[2][0][27] ,
         \s_mux2_signals[2][0][26] , \s_mux2_signals[2][0][25] ,
         \s_mux2_signals[2][0][24] , \s_mux2_signals[2][0][23] ,
         \s_mux2_signals[2][0][22] , \s_mux2_signals[2][0][21] ,
         \s_mux2_signals[2][0][20] , \s_mux2_signals[2][0][19] ,
         \s_mux2_signals[2][0][18] , \s_mux2_signals[2][0][17] ,
         \s_mux2_signals[2][0][16] , \s_mux2_signals[2][0][15] ,
         \s_mux2_signals[2][0][14] , \s_mux2_signals[2][0][13] ,
         \s_mux2_signals[2][0][12] , \s_mux2_signals[2][0][11] ,
         \s_mux2_signals[2][0][10] , \s_mux2_signals[2][0][9] ,
         \s_mux2_signals[2][0][8] , \s_mux2_signals[2][0][7] ,
         \s_mux2_signals[2][0][6] , \s_mux2_signals[2][0][5] ,
         \s_mux2_signals[2][0][4] , \s_mux2_signals[2][0][3] ,
         \s_mux2_signals[2][0][2] , \s_mux2_signals[2][0][1] ,
         \s_mux2_signals[2][0][0] , \s_mux2_signals[2][4][31] ,
         \s_mux2_signals[2][4][30] , \s_mux2_signals[2][4][29] ,
         \s_mux2_signals[2][4][28] , \s_mux2_signals[2][4][27] ,
         \s_mux2_signals[2][4][26] , \s_mux2_signals[2][4][25] ,
         \s_mux2_signals[2][4][24] , \s_mux2_signals[2][4][23] ,
         \s_mux2_signals[2][4][22] , \s_mux2_signals[2][4][21] ,
         \s_mux2_signals[2][4][20] , \s_mux2_signals[2][4][19] ,
         \s_mux2_signals[2][4][18] , \s_mux2_signals[2][4][17] ,
         \s_mux2_signals[2][4][16] , \s_mux2_signals[2][4][15] ,
         \s_mux2_signals[2][4][14] , \s_mux2_signals[2][4][13] ,
         \s_mux2_signals[2][4][12] , \s_mux2_signals[2][4][11] ,
         \s_mux2_signals[2][4][10] , \s_mux2_signals[2][4][9] ,
         \s_mux2_signals[2][4][8] , \s_mux2_signals[2][4][7] ,
         \s_mux2_signals[2][4][6] , \s_mux2_signals[2][4][5] ,
         \s_mux2_signals[2][4][4] , \s_mux2_signals[2][4][3] ,
         \s_mux2_signals[2][4][2] , \s_mux2_signals[2][4][1] ,
         \s_mux2_signals[2][4][0] , \s_mux2_signals[2][8][31] ,
         \s_mux2_signals[2][8][30] , \s_mux2_signals[2][8][29] ,
         \s_mux2_signals[2][8][28] , \s_mux2_signals[2][8][27] ,
         \s_mux2_signals[2][8][26] , \s_mux2_signals[2][8][25] ,
         \s_mux2_signals[2][8][24] , \s_mux2_signals[2][8][23] ,
         \s_mux2_signals[2][8][22] , \s_mux2_signals[2][8][21] ,
         \s_mux2_signals[2][8][20] , \s_mux2_signals[2][8][19] ,
         \s_mux2_signals[2][8][18] , \s_mux2_signals[2][8][17] ,
         \s_mux2_signals[2][8][16] , \s_mux2_signals[2][8][15] ,
         \s_mux2_signals[2][8][14] , \s_mux2_signals[2][8][13] ,
         \s_mux2_signals[2][8][12] , \s_mux2_signals[2][8][11] ,
         \s_mux2_signals[2][8][10] , \s_mux2_signals[2][8][9] ,
         \s_mux2_signals[2][8][8] , \s_mux2_signals[2][8][7] ,
         \s_mux2_signals[2][8][6] , \s_mux2_signals[2][8][5] ,
         \s_mux2_signals[2][8][4] , \s_mux2_signals[2][8][3] ,
         \s_mux2_signals[2][8][2] , \s_mux2_signals[2][8][1] ,
         \s_mux2_signals[2][8][0] , \s_mux2_signals[2][12][31] ,
         \s_mux2_signals[2][12][30] , \s_mux2_signals[2][12][29] ,
         \s_mux2_signals[2][12][28] , \s_mux2_signals[2][12][27] ,
         \s_mux2_signals[2][12][26] , \s_mux2_signals[2][12][25] ,
         \s_mux2_signals[2][12][24] , \s_mux2_signals[2][12][23] ,
         \s_mux2_signals[2][12][22] , \s_mux2_signals[2][12][21] ,
         \s_mux2_signals[2][12][20] , \s_mux2_signals[2][12][19] ,
         \s_mux2_signals[2][12][18] , \s_mux2_signals[2][12][17] ,
         \s_mux2_signals[2][12][16] , \s_mux2_signals[2][12][15] ,
         \s_mux2_signals[2][12][14] , \s_mux2_signals[2][12][13] ,
         \s_mux2_signals[2][12][12] , \s_mux2_signals[2][12][11] ,
         \s_mux2_signals[2][12][10] , \s_mux2_signals[2][12][9] ,
         \s_mux2_signals[2][12][8] , \s_mux2_signals[2][12][7] ,
         \s_mux2_signals[2][12][6] , \s_mux2_signals[2][12][5] ,
         \s_mux2_signals[2][12][4] , \s_mux2_signals[2][12][3] ,
         \s_mux2_signals[2][12][2] , \s_mux2_signals[2][12][1] ,
         \s_mux2_signals[2][12][0] , \s_mux2_signals[2][16][31] ,
         \s_mux2_signals[2][16][30] , \s_mux2_signals[2][16][29] ,
         \s_mux2_signals[2][16][28] , \s_mux2_signals[2][16][27] ,
         \s_mux2_signals[2][16][26] , \s_mux2_signals[2][16][25] ,
         \s_mux2_signals[2][16][24] , \s_mux2_signals[2][16][23] ,
         \s_mux2_signals[2][16][22] , \s_mux2_signals[2][16][21] ,
         \s_mux2_signals[2][16][20] , \s_mux2_signals[2][16][19] ,
         \s_mux2_signals[2][16][18] , \s_mux2_signals[2][16][17] ,
         \s_mux2_signals[2][16][16] , \s_mux2_signals[2][16][15] ,
         \s_mux2_signals[2][16][14] , \s_mux2_signals[2][16][13] ,
         \s_mux2_signals[2][16][12] , \s_mux2_signals[2][16][11] ,
         \s_mux2_signals[2][16][10] , \s_mux2_signals[2][16][9] ,
         \s_mux2_signals[2][16][8] , \s_mux2_signals[2][16][7] ,
         \s_mux2_signals[2][16][6] , \s_mux2_signals[2][16][5] ,
         \s_mux2_signals[2][16][4] , \s_mux2_signals[2][16][3] ,
         \s_mux2_signals[2][16][2] , \s_mux2_signals[2][16][1] ,
         \s_mux2_signals[2][16][0] , \s_mux2_signals[2][20][31] ,
         \s_mux2_signals[2][20][30] , \s_mux2_signals[2][20][29] ,
         \s_mux2_signals[2][20][28] , \s_mux2_signals[2][20][27] ,
         \s_mux2_signals[2][20][26] , \s_mux2_signals[2][20][25] ,
         \s_mux2_signals[2][20][24] , \s_mux2_signals[2][20][23] ,
         \s_mux2_signals[2][20][22] , \s_mux2_signals[2][20][21] ,
         \s_mux2_signals[2][20][20] , \s_mux2_signals[2][20][19] ,
         \s_mux2_signals[2][20][18] , \s_mux2_signals[2][20][17] ,
         \s_mux2_signals[2][20][16] , \s_mux2_signals[2][20][15] ,
         \s_mux2_signals[2][20][14] , \s_mux2_signals[2][20][13] ,
         \s_mux2_signals[2][20][12] , \s_mux2_signals[2][20][11] ,
         \s_mux2_signals[2][20][10] , \s_mux2_signals[2][20][9] ,
         \s_mux2_signals[2][20][8] , \s_mux2_signals[2][20][7] ,
         \s_mux2_signals[2][20][6] , \s_mux2_signals[2][20][5] ,
         \s_mux2_signals[2][20][4] , \s_mux2_signals[2][20][3] ,
         \s_mux2_signals[2][20][2] , \s_mux2_signals[2][20][1] ,
         \s_mux2_signals[2][20][0] , \s_mux2_signals[2][24][31] ,
         \s_mux2_signals[2][24][30] , \s_mux2_signals[2][24][29] ,
         \s_mux2_signals[2][24][28] , \s_mux2_signals[2][24][27] ,
         \s_mux2_signals[2][24][26] , \s_mux2_signals[2][24][25] ,
         \s_mux2_signals[2][24][24] , \s_mux2_signals[2][24][23] ,
         \s_mux2_signals[2][24][22] , \s_mux2_signals[2][24][21] ,
         \s_mux2_signals[2][24][20] , \s_mux2_signals[2][24][19] ,
         \s_mux2_signals[2][24][18] , \s_mux2_signals[2][24][17] ,
         \s_mux2_signals[2][24][16] , \s_mux2_signals[2][24][15] ,
         \s_mux2_signals[2][24][14] , \s_mux2_signals[2][24][13] ,
         \s_mux2_signals[2][24][12] , \s_mux2_signals[2][24][11] ,
         \s_mux2_signals[2][24][10] , \s_mux2_signals[2][24][9] ,
         \s_mux2_signals[2][24][8] , \s_mux2_signals[2][24][7] ,
         \s_mux2_signals[2][24][6] , \s_mux2_signals[2][24][5] ,
         \s_mux2_signals[2][24][4] , \s_mux2_signals[2][24][3] ,
         \s_mux2_signals[2][24][2] , \s_mux2_signals[2][24][1] ,
         \s_mux2_signals[2][24][0] , \s_mux2_signals[2][28][31] ,
         \s_mux2_signals[2][28][30] , \s_mux2_signals[2][28][29] ,
         \s_mux2_signals[2][28][28] , \s_mux2_signals[2][28][27] ,
         \s_mux2_signals[2][28][26] , \s_mux2_signals[2][28][25] ,
         \s_mux2_signals[2][28][24] , \s_mux2_signals[2][28][23] ,
         \s_mux2_signals[2][28][22] , \s_mux2_signals[2][28][21] ,
         \s_mux2_signals[2][28][20] , \s_mux2_signals[2][28][19] ,
         \s_mux2_signals[2][28][18] , \s_mux2_signals[2][28][17] ,
         \s_mux2_signals[2][28][16] , \s_mux2_signals[2][28][15] ,
         \s_mux2_signals[2][28][14] , \s_mux2_signals[2][28][13] ,
         \s_mux2_signals[2][28][12] , \s_mux2_signals[2][28][11] ,
         \s_mux2_signals[2][28][10] , \s_mux2_signals[2][28][9] ,
         \s_mux2_signals[2][28][8] , \s_mux2_signals[2][28][7] ,
         \s_mux2_signals[2][28][6] , \s_mux2_signals[2][28][5] ,
         \s_mux2_signals[2][28][4] , \s_mux2_signals[2][28][3] ,
         \s_mux2_signals[2][28][2] , \s_mux2_signals[2][28][1] ,
         \s_mux2_signals[2][28][0] , \s_mux2_signals[3][0][31] ,
         \s_mux2_signals[3][0][30] , \s_mux2_signals[3][0][29] ,
         \s_mux2_signals[3][0][28] , \s_mux2_signals[3][0][27] ,
         \s_mux2_signals[3][0][26] , \s_mux2_signals[3][0][25] ,
         \s_mux2_signals[3][0][24] , \s_mux2_signals[3][0][23] ,
         \s_mux2_signals[3][0][22] , \s_mux2_signals[3][0][21] ,
         \s_mux2_signals[3][0][20] , \s_mux2_signals[3][0][19] ,
         \s_mux2_signals[3][0][18] , \s_mux2_signals[3][0][17] ,
         \s_mux2_signals[3][0][16] , \s_mux2_signals[3][0][15] ,
         \s_mux2_signals[3][0][14] , \s_mux2_signals[3][0][13] ,
         \s_mux2_signals[3][0][12] , \s_mux2_signals[3][0][11] ,
         \s_mux2_signals[3][0][10] , \s_mux2_signals[3][0][9] ,
         \s_mux2_signals[3][0][8] , \s_mux2_signals[3][0][7] ,
         \s_mux2_signals[3][0][6] , \s_mux2_signals[3][0][5] ,
         \s_mux2_signals[3][0][4] , \s_mux2_signals[3][0][3] ,
         \s_mux2_signals[3][0][2] , \s_mux2_signals[3][0][1] ,
         \s_mux2_signals[3][0][0] , \s_mux2_signals[3][8][31] ,
         \s_mux2_signals[3][8][30] , \s_mux2_signals[3][8][29] ,
         \s_mux2_signals[3][8][28] , \s_mux2_signals[3][8][27] ,
         \s_mux2_signals[3][8][26] , \s_mux2_signals[3][8][25] ,
         \s_mux2_signals[3][8][24] , \s_mux2_signals[3][8][23] ,
         \s_mux2_signals[3][8][22] , \s_mux2_signals[3][8][21] ,
         \s_mux2_signals[3][8][20] , \s_mux2_signals[3][8][19] ,
         \s_mux2_signals[3][8][18] , \s_mux2_signals[3][8][17] ,
         \s_mux2_signals[3][8][16] , \s_mux2_signals[3][8][15] ,
         \s_mux2_signals[3][8][14] , \s_mux2_signals[3][8][13] ,
         \s_mux2_signals[3][8][12] , \s_mux2_signals[3][8][11] ,
         \s_mux2_signals[3][8][10] , \s_mux2_signals[3][8][9] ,
         \s_mux2_signals[3][8][8] , \s_mux2_signals[3][8][7] ,
         \s_mux2_signals[3][8][6] , \s_mux2_signals[3][8][5] ,
         \s_mux2_signals[3][8][4] , \s_mux2_signals[3][8][3] ,
         \s_mux2_signals[3][8][2] , \s_mux2_signals[3][8][1] ,
         \s_mux2_signals[3][8][0] , \s_mux2_signals[3][16][31] ,
         \s_mux2_signals[3][16][30] , \s_mux2_signals[3][16][29] ,
         \s_mux2_signals[3][16][28] , \s_mux2_signals[3][16][27] ,
         \s_mux2_signals[3][16][26] , \s_mux2_signals[3][16][25] ,
         \s_mux2_signals[3][16][24] , \s_mux2_signals[3][16][23] ,
         \s_mux2_signals[3][16][22] , \s_mux2_signals[3][16][21] ,
         \s_mux2_signals[3][16][20] , \s_mux2_signals[3][16][19] ,
         \s_mux2_signals[3][16][18] , \s_mux2_signals[3][16][17] ,
         \s_mux2_signals[3][16][16] , \s_mux2_signals[3][16][15] ,
         \s_mux2_signals[3][16][14] , \s_mux2_signals[3][16][13] ,
         \s_mux2_signals[3][16][12] , \s_mux2_signals[3][16][11] ,
         \s_mux2_signals[3][16][10] , \s_mux2_signals[3][16][9] ,
         \s_mux2_signals[3][16][8] , \s_mux2_signals[3][16][7] ,
         \s_mux2_signals[3][16][6] , \s_mux2_signals[3][16][5] ,
         \s_mux2_signals[3][16][4] , \s_mux2_signals[3][16][3] ,
         \s_mux2_signals[3][16][2] , \s_mux2_signals[3][16][1] ,
         \s_mux2_signals[3][16][0] , \s_mux2_signals[3][24][31] ,
         \s_mux2_signals[3][24][30] , \s_mux2_signals[3][24][29] ,
         \s_mux2_signals[3][24][28] , \s_mux2_signals[3][24][27] ,
         \s_mux2_signals[3][24][26] , \s_mux2_signals[3][24][25] ,
         \s_mux2_signals[3][24][24] , \s_mux2_signals[3][24][23] ,
         \s_mux2_signals[3][24][22] , \s_mux2_signals[3][24][21] ,
         \s_mux2_signals[3][24][20] , \s_mux2_signals[3][24][19] ,
         \s_mux2_signals[3][24][18] , \s_mux2_signals[3][24][17] ,
         \s_mux2_signals[3][24][16] , \s_mux2_signals[3][24][15] ,
         \s_mux2_signals[3][24][14] , \s_mux2_signals[3][24][13] ,
         \s_mux2_signals[3][24][12] , \s_mux2_signals[3][24][11] ,
         \s_mux2_signals[3][24][10] , \s_mux2_signals[3][24][9] ,
         \s_mux2_signals[3][24][8] , \s_mux2_signals[3][24][7] ,
         \s_mux2_signals[3][24][6] , \s_mux2_signals[3][24][5] ,
         \s_mux2_signals[3][24][4] , \s_mux2_signals[3][24][3] ,
         \s_mux2_signals[3][24][2] , \s_mux2_signals[3][24][1] ,
         \s_mux2_signals[3][24][0] , \s_mux2_signals[4][0][31] ,
         \s_mux2_signals[4][0][30] , \s_mux2_signals[4][0][29] ,
         \s_mux2_signals[4][0][28] , \s_mux2_signals[4][0][27] ,
         \s_mux2_signals[4][0][26] , \s_mux2_signals[4][0][25] ,
         \s_mux2_signals[4][0][24] , \s_mux2_signals[4][0][23] ,
         \s_mux2_signals[4][0][22] , \s_mux2_signals[4][0][21] ,
         \s_mux2_signals[4][0][20] , \s_mux2_signals[4][0][19] ,
         \s_mux2_signals[4][0][18] , \s_mux2_signals[4][0][17] ,
         \s_mux2_signals[4][0][16] , \s_mux2_signals[4][0][15] ,
         \s_mux2_signals[4][0][14] , \s_mux2_signals[4][0][13] ,
         \s_mux2_signals[4][0][12] , \s_mux2_signals[4][0][11] ,
         \s_mux2_signals[4][0][10] , \s_mux2_signals[4][0][9] ,
         \s_mux2_signals[4][0][8] , \s_mux2_signals[4][0][7] ,
         \s_mux2_signals[4][0][6] , \s_mux2_signals[4][0][5] ,
         \s_mux2_signals[4][0][4] , \s_mux2_signals[4][0][3] ,
         \s_mux2_signals[4][0][2] , \s_mux2_signals[4][0][1] ,
         \s_mux2_signals[4][0][0] , \s_mux2_signals[4][16][31] ,
         \s_mux2_signals[4][16][30] , \s_mux2_signals[4][16][29] ,
         \s_mux2_signals[4][16][28] , \s_mux2_signals[4][16][27] ,
         \s_mux2_signals[4][16][26] , \s_mux2_signals[4][16][25] ,
         \s_mux2_signals[4][16][24] , \s_mux2_signals[4][16][23] ,
         \s_mux2_signals[4][16][22] , \s_mux2_signals[4][16][21] ,
         \s_mux2_signals[4][16][20] , \s_mux2_signals[4][16][19] ,
         \s_mux2_signals[4][16][18] , \s_mux2_signals[4][16][17] ,
         \s_mux2_signals[4][16][16] , \s_mux2_signals[4][16][15] ,
         \s_mux2_signals[4][16][14] , \s_mux2_signals[4][16][13] ,
         \s_mux2_signals[4][16][12] , \s_mux2_signals[4][16][11] ,
         \s_mux2_signals[4][16][10] , \s_mux2_signals[4][16][9] ,
         \s_mux2_signals[4][16][8] , \s_mux2_signals[4][16][7] ,
         \s_mux2_signals[4][16][6] , \s_mux2_signals[4][16][5] ,
         \s_mux2_signals[4][16][4] , \s_mux2_signals[4][16][3] ,
         \s_mux2_signals[4][16][2] , \s_mux2_signals[4][16][1] ,
         \s_mux2_signals[4][16][0] , \s_mux1_signals[1][0][31] ,
         \s_mux1_signals[1][0][30] , \s_mux1_signals[1][0][29] ,
         \s_mux1_signals[1][0][28] , \s_mux1_signals[1][0][27] ,
         \s_mux1_signals[1][0][26] , \s_mux1_signals[1][0][25] ,
         \s_mux1_signals[1][0][24] , \s_mux1_signals[1][0][23] ,
         \s_mux1_signals[1][0][22] , \s_mux1_signals[1][0][21] ,
         \s_mux1_signals[1][0][20] , \s_mux1_signals[1][0][19] ,
         \s_mux1_signals[1][0][18] , \s_mux1_signals[1][0][17] ,
         \s_mux1_signals[1][0][16] , \s_mux1_signals[1][0][15] ,
         \s_mux1_signals[1][0][14] , \s_mux1_signals[1][0][13] ,
         \s_mux1_signals[1][0][12] , \s_mux1_signals[1][0][11] ,
         \s_mux1_signals[1][0][10] , \s_mux1_signals[1][0][9] ,
         \s_mux1_signals[1][0][8] , \s_mux1_signals[1][0][7] ,
         \s_mux1_signals[1][0][6] , \s_mux1_signals[1][0][5] ,
         \s_mux1_signals[1][0][4] , \s_mux1_signals[1][0][3] ,
         \s_mux1_signals[1][0][2] , \s_mux1_signals[1][0][1] ,
         \s_mux1_signals[1][0][0] , \s_mux1_signals[1][2][31] ,
         \s_mux1_signals[1][2][30] , \s_mux1_signals[1][2][29] ,
         \s_mux1_signals[1][2][28] , \s_mux1_signals[1][2][27] ,
         \s_mux1_signals[1][2][26] , \s_mux1_signals[1][2][25] ,
         \s_mux1_signals[1][2][24] , \s_mux1_signals[1][2][23] ,
         \s_mux1_signals[1][2][22] , \s_mux1_signals[1][2][21] ,
         \s_mux1_signals[1][2][20] , \s_mux1_signals[1][2][19] ,
         \s_mux1_signals[1][2][18] , \s_mux1_signals[1][2][17] ,
         \s_mux1_signals[1][2][16] , \s_mux1_signals[1][2][15] ,
         \s_mux1_signals[1][2][14] , \s_mux1_signals[1][2][13] ,
         \s_mux1_signals[1][2][12] , \s_mux1_signals[1][2][11] ,
         \s_mux1_signals[1][2][10] , \s_mux1_signals[1][2][9] ,
         \s_mux1_signals[1][2][8] , \s_mux1_signals[1][2][7] ,
         \s_mux1_signals[1][2][6] , \s_mux1_signals[1][2][5] ,
         \s_mux1_signals[1][2][4] , \s_mux1_signals[1][2][3] ,
         \s_mux1_signals[1][2][2] , \s_mux1_signals[1][2][1] ,
         \s_mux1_signals[1][2][0] , \s_mux1_signals[1][4][31] ,
         \s_mux1_signals[1][4][30] , \s_mux1_signals[1][4][29] ,
         \s_mux1_signals[1][4][28] , \s_mux1_signals[1][4][27] ,
         \s_mux1_signals[1][4][26] , \s_mux1_signals[1][4][25] ,
         \s_mux1_signals[1][4][24] , \s_mux1_signals[1][4][23] ,
         \s_mux1_signals[1][4][22] , \s_mux1_signals[1][4][21] ,
         \s_mux1_signals[1][4][20] , \s_mux1_signals[1][4][19] ,
         \s_mux1_signals[1][4][18] , \s_mux1_signals[1][4][17] ,
         \s_mux1_signals[1][4][16] , \s_mux1_signals[1][4][15] ,
         \s_mux1_signals[1][4][14] , \s_mux1_signals[1][4][13] ,
         \s_mux1_signals[1][4][12] , \s_mux1_signals[1][4][11] ,
         \s_mux1_signals[1][4][10] , \s_mux1_signals[1][4][9] ,
         \s_mux1_signals[1][4][8] , \s_mux1_signals[1][4][7] ,
         \s_mux1_signals[1][4][6] , \s_mux1_signals[1][4][5] ,
         \s_mux1_signals[1][4][4] , \s_mux1_signals[1][4][3] ,
         \s_mux1_signals[1][4][2] , \s_mux1_signals[1][4][1] ,
         \s_mux1_signals[1][4][0] , \s_mux1_signals[1][6][31] ,
         \s_mux1_signals[1][6][30] , \s_mux1_signals[1][6][29] ,
         \s_mux1_signals[1][6][28] , \s_mux1_signals[1][6][27] ,
         \s_mux1_signals[1][6][26] , \s_mux1_signals[1][6][25] ,
         \s_mux1_signals[1][6][24] , \s_mux1_signals[1][6][23] ,
         \s_mux1_signals[1][6][22] , \s_mux1_signals[1][6][21] ,
         \s_mux1_signals[1][6][20] , \s_mux1_signals[1][6][19] ,
         \s_mux1_signals[1][6][18] , \s_mux1_signals[1][6][17] ,
         \s_mux1_signals[1][6][16] , \s_mux1_signals[1][6][15] ,
         \s_mux1_signals[1][6][14] , \s_mux1_signals[1][6][13] ,
         \s_mux1_signals[1][6][12] , \s_mux1_signals[1][6][11] ,
         \s_mux1_signals[1][6][10] , \s_mux1_signals[1][6][9] ,
         \s_mux1_signals[1][6][8] , \s_mux1_signals[1][6][7] ,
         \s_mux1_signals[1][6][6] , \s_mux1_signals[1][6][5] ,
         \s_mux1_signals[1][6][4] , \s_mux1_signals[1][6][3] ,
         \s_mux1_signals[1][6][2] , \s_mux1_signals[1][6][1] ,
         \s_mux1_signals[1][6][0] , \s_mux1_signals[1][8][31] ,
         \s_mux1_signals[1][8][30] , \s_mux1_signals[1][8][29] ,
         \s_mux1_signals[1][8][28] , \s_mux1_signals[1][8][27] ,
         \s_mux1_signals[1][8][26] , \s_mux1_signals[1][8][25] ,
         \s_mux1_signals[1][8][24] , \s_mux1_signals[1][8][23] ,
         \s_mux1_signals[1][8][22] , \s_mux1_signals[1][8][21] ,
         \s_mux1_signals[1][8][20] , \s_mux1_signals[1][8][19] ,
         \s_mux1_signals[1][8][18] , \s_mux1_signals[1][8][17] ,
         \s_mux1_signals[1][8][16] , \s_mux1_signals[1][8][15] ,
         \s_mux1_signals[1][8][14] , \s_mux1_signals[1][8][13] ,
         \s_mux1_signals[1][8][12] , \s_mux1_signals[1][8][11] ,
         \s_mux1_signals[1][8][10] , \s_mux1_signals[1][8][9] ,
         \s_mux1_signals[1][8][8] , \s_mux1_signals[1][8][7] ,
         \s_mux1_signals[1][8][6] , \s_mux1_signals[1][8][5] ,
         \s_mux1_signals[1][8][4] , \s_mux1_signals[1][8][3] ,
         \s_mux1_signals[1][8][2] , \s_mux1_signals[1][8][1] ,
         \s_mux1_signals[1][8][0] , \s_mux1_signals[1][10][31] ,
         \s_mux1_signals[1][10][30] , \s_mux1_signals[1][10][29] ,
         \s_mux1_signals[1][10][28] , \s_mux1_signals[1][10][27] ,
         \s_mux1_signals[1][10][26] , \s_mux1_signals[1][10][25] ,
         \s_mux1_signals[1][10][24] , \s_mux1_signals[1][10][23] ,
         \s_mux1_signals[1][10][22] , \s_mux1_signals[1][10][21] ,
         \s_mux1_signals[1][10][20] , \s_mux1_signals[1][10][19] ,
         \s_mux1_signals[1][10][18] , \s_mux1_signals[1][10][17] ,
         \s_mux1_signals[1][10][16] , \s_mux1_signals[1][10][15] ,
         \s_mux1_signals[1][10][14] , \s_mux1_signals[1][10][13] ,
         \s_mux1_signals[1][10][12] , \s_mux1_signals[1][10][11] ,
         \s_mux1_signals[1][10][10] , \s_mux1_signals[1][10][9] ,
         \s_mux1_signals[1][10][8] , \s_mux1_signals[1][10][7] ,
         \s_mux1_signals[1][10][6] , \s_mux1_signals[1][10][5] ,
         \s_mux1_signals[1][10][4] , \s_mux1_signals[1][10][3] ,
         \s_mux1_signals[1][10][2] , \s_mux1_signals[1][10][1] ,
         \s_mux1_signals[1][10][0] , \s_mux1_signals[1][12][31] ,
         \s_mux1_signals[1][12][30] , \s_mux1_signals[1][12][29] ,
         \s_mux1_signals[1][12][28] , \s_mux1_signals[1][12][27] ,
         \s_mux1_signals[1][12][26] , \s_mux1_signals[1][12][25] ,
         \s_mux1_signals[1][12][24] , \s_mux1_signals[1][12][23] ,
         \s_mux1_signals[1][12][22] , \s_mux1_signals[1][12][21] ,
         \s_mux1_signals[1][12][20] , \s_mux1_signals[1][12][19] ,
         \s_mux1_signals[1][12][18] , \s_mux1_signals[1][12][17] ,
         \s_mux1_signals[1][12][16] , \s_mux1_signals[1][12][15] ,
         \s_mux1_signals[1][12][14] , \s_mux1_signals[1][12][13] ,
         \s_mux1_signals[1][12][12] , \s_mux1_signals[1][12][11] ,
         \s_mux1_signals[1][12][10] , \s_mux1_signals[1][12][9] ,
         \s_mux1_signals[1][12][8] , \s_mux1_signals[1][12][7] ,
         \s_mux1_signals[1][12][6] , \s_mux1_signals[1][12][5] ,
         \s_mux1_signals[1][12][4] , \s_mux1_signals[1][12][3] ,
         \s_mux1_signals[1][12][2] , \s_mux1_signals[1][12][1] ,
         \s_mux1_signals[1][12][0] , \s_mux1_signals[1][14][31] ,
         \s_mux1_signals[1][14][30] , \s_mux1_signals[1][14][29] ,
         \s_mux1_signals[1][14][28] , \s_mux1_signals[1][14][27] ,
         \s_mux1_signals[1][14][26] , \s_mux1_signals[1][14][25] ,
         \s_mux1_signals[1][14][24] , \s_mux1_signals[1][14][23] ,
         \s_mux1_signals[1][14][22] , \s_mux1_signals[1][14][21] ,
         \s_mux1_signals[1][14][20] , \s_mux1_signals[1][14][19] ,
         \s_mux1_signals[1][14][18] , \s_mux1_signals[1][14][17] ,
         \s_mux1_signals[1][14][16] , \s_mux1_signals[1][14][15] ,
         \s_mux1_signals[1][14][14] , \s_mux1_signals[1][14][13] ,
         \s_mux1_signals[1][14][12] , \s_mux1_signals[1][14][11] ,
         \s_mux1_signals[1][14][10] , \s_mux1_signals[1][14][9] ,
         \s_mux1_signals[1][14][8] , \s_mux1_signals[1][14][7] ,
         \s_mux1_signals[1][14][6] , \s_mux1_signals[1][14][5] ,
         \s_mux1_signals[1][14][4] , \s_mux1_signals[1][14][3] ,
         \s_mux1_signals[1][14][2] , \s_mux1_signals[1][14][1] ,
         \s_mux1_signals[1][14][0] , \s_mux1_signals[1][16][31] ,
         \s_mux1_signals[1][16][30] , \s_mux1_signals[1][16][29] ,
         \s_mux1_signals[1][16][28] , \s_mux1_signals[1][16][27] ,
         \s_mux1_signals[1][16][26] , \s_mux1_signals[1][16][25] ,
         \s_mux1_signals[1][16][24] , \s_mux1_signals[1][16][23] ,
         \s_mux1_signals[1][16][22] , \s_mux1_signals[1][16][21] ,
         \s_mux1_signals[1][16][20] , \s_mux1_signals[1][16][19] ,
         \s_mux1_signals[1][16][18] , \s_mux1_signals[1][16][17] ,
         \s_mux1_signals[1][16][16] , \s_mux1_signals[1][16][15] ,
         \s_mux1_signals[1][16][14] , \s_mux1_signals[1][16][13] ,
         \s_mux1_signals[1][16][12] , \s_mux1_signals[1][16][11] ,
         \s_mux1_signals[1][16][10] , \s_mux1_signals[1][16][9] ,
         \s_mux1_signals[1][16][8] , \s_mux1_signals[1][16][7] ,
         \s_mux1_signals[1][16][6] , \s_mux1_signals[1][16][5] ,
         \s_mux1_signals[1][16][4] , \s_mux1_signals[1][16][3] ,
         \s_mux1_signals[1][16][2] , \s_mux1_signals[1][16][1] ,
         \s_mux1_signals[1][16][0] , \s_mux1_signals[1][18][31] ,
         \s_mux1_signals[1][18][30] , \s_mux1_signals[1][18][29] ,
         \s_mux1_signals[1][18][28] , \s_mux1_signals[1][18][27] ,
         \s_mux1_signals[1][18][26] , \s_mux1_signals[1][18][25] ,
         \s_mux1_signals[1][18][24] , \s_mux1_signals[1][18][23] ,
         \s_mux1_signals[1][18][22] , \s_mux1_signals[1][18][21] ,
         \s_mux1_signals[1][18][20] , \s_mux1_signals[1][18][19] ,
         \s_mux1_signals[1][18][18] , \s_mux1_signals[1][18][17] ,
         \s_mux1_signals[1][18][16] , \s_mux1_signals[1][18][15] ,
         \s_mux1_signals[1][18][14] , \s_mux1_signals[1][18][13] ,
         \s_mux1_signals[1][18][12] , \s_mux1_signals[1][18][11] ,
         \s_mux1_signals[1][18][10] , \s_mux1_signals[1][18][9] ,
         \s_mux1_signals[1][18][8] , \s_mux1_signals[1][18][7] ,
         \s_mux1_signals[1][18][6] , \s_mux1_signals[1][18][5] ,
         \s_mux1_signals[1][18][4] , \s_mux1_signals[1][18][3] ,
         \s_mux1_signals[1][18][2] , \s_mux1_signals[1][18][1] ,
         \s_mux1_signals[1][18][0] , \s_mux1_signals[1][20][31] ,
         \s_mux1_signals[1][20][30] , \s_mux1_signals[1][20][29] ,
         \s_mux1_signals[1][20][28] , \s_mux1_signals[1][20][27] ,
         \s_mux1_signals[1][20][26] , \s_mux1_signals[1][20][25] ,
         \s_mux1_signals[1][20][24] , \s_mux1_signals[1][20][23] ,
         \s_mux1_signals[1][20][22] , \s_mux1_signals[1][20][21] ,
         \s_mux1_signals[1][20][20] , \s_mux1_signals[1][20][19] ,
         \s_mux1_signals[1][20][18] , \s_mux1_signals[1][20][17] ,
         \s_mux1_signals[1][20][16] , \s_mux1_signals[1][20][15] ,
         \s_mux1_signals[1][20][14] , \s_mux1_signals[1][20][13] ,
         \s_mux1_signals[1][20][12] , \s_mux1_signals[1][20][11] ,
         \s_mux1_signals[1][20][10] , \s_mux1_signals[1][20][9] ,
         \s_mux1_signals[1][20][8] , \s_mux1_signals[1][20][7] ,
         \s_mux1_signals[1][20][6] , \s_mux1_signals[1][20][5] ,
         \s_mux1_signals[1][20][4] , \s_mux1_signals[1][20][3] ,
         \s_mux1_signals[1][20][2] , \s_mux1_signals[1][20][1] ,
         \s_mux1_signals[1][20][0] , \s_mux1_signals[1][22][31] ,
         \s_mux1_signals[1][22][30] , \s_mux1_signals[1][22][29] ,
         \s_mux1_signals[1][22][28] , \s_mux1_signals[1][22][27] ,
         \s_mux1_signals[1][22][26] , \s_mux1_signals[1][22][25] ,
         \s_mux1_signals[1][22][24] , \s_mux1_signals[1][22][23] ,
         \s_mux1_signals[1][22][22] , \s_mux1_signals[1][22][21] ,
         \s_mux1_signals[1][22][20] , \s_mux1_signals[1][22][19] ,
         \s_mux1_signals[1][22][18] , \s_mux1_signals[1][22][17] ,
         \s_mux1_signals[1][22][16] , \s_mux1_signals[1][22][15] ,
         \s_mux1_signals[1][22][14] , \s_mux1_signals[1][22][13] ,
         \s_mux1_signals[1][22][12] , \s_mux1_signals[1][22][11] ,
         \s_mux1_signals[1][22][10] , \s_mux1_signals[1][22][9] ,
         \s_mux1_signals[1][22][8] , \s_mux1_signals[1][22][7] ,
         \s_mux1_signals[1][22][6] , \s_mux1_signals[1][22][5] ,
         \s_mux1_signals[1][22][4] , \s_mux1_signals[1][22][3] ,
         \s_mux1_signals[1][22][2] , \s_mux1_signals[1][22][1] ,
         \s_mux1_signals[1][22][0] , \s_mux1_signals[1][24][31] ,
         \s_mux1_signals[1][24][30] , \s_mux1_signals[1][24][29] ,
         \s_mux1_signals[1][24][28] , \s_mux1_signals[1][24][27] ,
         \s_mux1_signals[1][24][26] , \s_mux1_signals[1][24][25] ,
         \s_mux1_signals[1][24][24] , \s_mux1_signals[1][24][23] ,
         \s_mux1_signals[1][24][22] , \s_mux1_signals[1][24][21] ,
         \s_mux1_signals[1][24][20] , \s_mux1_signals[1][24][19] ,
         \s_mux1_signals[1][24][18] , \s_mux1_signals[1][24][17] ,
         \s_mux1_signals[1][24][16] , \s_mux1_signals[1][24][15] ,
         \s_mux1_signals[1][24][14] , \s_mux1_signals[1][24][13] ,
         \s_mux1_signals[1][24][12] , \s_mux1_signals[1][24][11] ,
         \s_mux1_signals[1][24][10] , \s_mux1_signals[1][24][9] ,
         \s_mux1_signals[1][24][8] , \s_mux1_signals[1][24][7] ,
         \s_mux1_signals[1][24][6] , \s_mux1_signals[1][24][5] ,
         \s_mux1_signals[1][24][4] , \s_mux1_signals[1][24][3] ,
         \s_mux1_signals[1][24][2] , \s_mux1_signals[1][24][1] ,
         \s_mux1_signals[1][24][0] , \s_mux1_signals[1][26][31] ,
         \s_mux1_signals[1][26][30] , \s_mux1_signals[1][26][29] ,
         \s_mux1_signals[1][26][28] , \s_mux1_signals[1][26][27] ,
         \s_mux1_signals[1][26][26] , \s_mux1_signals[1][26][25] ,
         \s_mux1_signals[1][26][24] , \s_mux1_signals[1][26][23] ,
         \s_mux1_signals[1][26][22] , \s_mux1_signals[1][26][21] ,
         \s_mux1_signals[1][26][20] , \s_mux1_signals[1][26][19] ,
         \s_mux1_signals[1][26][18] , \s_mux1_signals[1][26][17] ,
         \s_mux1_signals[1][26][16] , \s_mux1_signals[1][26][15] ,
         \s_mux1_signals[1][26][14] , \s_mux1_signals[1][26][13] ,
         \s_mux1_signals[1][26][12] , \s_mux1_signals[1][26][11] ,
         \s_mux1_signals[1][26][10] , \s_mux1_signals[1][26][9] ,
         \s_mux1_signals[1][26][8] , \s_mux1_signals[1][26][7] ,
         \s_mux1_signals[1][26][6] , \s_mux1_signals[1][26][5] ,
         \s_mux1_signals[1][26][4] , \s_mux1_signals[1][26][3] ,
         \s_mux1_signals[1][26][2] , \s_mux1_signals[1][26][1] ,
         \s_mux1_signals[1][26][0] , \s_mux1_signals[1][28][31] ,
         \s_mux1_signals[1][28][30] , \s_mux1_signals[1][28][29] ,
         \s_mux1_signals[1][28][28] , \s_mux1_signals[1][28][27] ,
         \s_mux1_signals[1][28][26] , \s_mux1_signals[1][28][25] ,
         \s_mux1_signals[1][28][24] , \s_mux1_signals[1][28][23] ,
         \s_mux1_signals[1][28][22] , \s_mux1_signals[1][28][21] ,
         \s_mux1_signals[1][28][20] , \s_mux1_signals[1][28][19] ,
         \s_mux1_signals[1][28][18] , \s_mux1_signals[1][28][17] ,
         \s_mux1_signals[1][28][16] , \s_mux1_signals[1][28][15] ,
         \s_mux1_signals[1][28][14] , \s_mux1_signals[1][28][13] ,
         \s_mux1_signals[1][28][12] , \s_mux1_signals[1][28][11] ,
         \s_mux1_signals[1][28][10] , \s_mux1_signals[1][28][9] ,
         \s_mux1_signals[1][28][8] , \s_mux1_signals[1][28][7] ,
         \s_mux1_signals[1][28][6] , \s_mux1_signals[1][28][5] ,
         \s_mux1_signals[1][28][4] , \s_mux1_signals[1][28][3] ,
         \s_mux1_signals[1][28][2] , \s_mux1_signals[1][28][1] ,
         \s_mux1_signals[1][28][0] , \s_mux1_signals[1][30][31] ,
         \s_mux1_signals[1][30][30] , \s_mux1_signals[1][30][29] ,
         \s_mux1_signals[1][30][28] , \s_mux1_signals[1][30][27] ,
         \s_mux1_signals[1][30][26] , \s_mux1_signals[1][30][25] ,
         \s_mux1_signals[1][30][24] , \s_mux1_signals[1][30][23] ,
         \s_mux1_signals[1][30][22] , \s_mux1_signals[1][30][21] ,
         \s_mux1_signals[1][30][20] , \s_mux1_signals[1][30][19] ,
         \s_mux1_signals[1][30][18] , \s_mux1_signals[1][30][17] ,
         \s_mux1_signals[1][30][16] , \s_mux1_signals[1][30][15] ,
         \s_mux1_signals[1][30][14] , \s_mux1_signals[1][30][13] ,
         \s_mux1_signals[1][30][12] , \s_mux1_signals[1][30][11] ,
         \s_mux1_signals[1][30][10] , \s_mux1_signals[1][30][9] ,
         \s_mux1_signals[1][30][8] , \s_mux1_signals[1][30][7] ,
         \s_mux1_signals[1][30][6] , \s_mux1_signals[1][30][5] ,
         \s_mux1_signals[1][30][4] , \s_mux1_signals[1][30][3] ,
         \s_mux1_signals[1][30][2] , \s_mux1_signals[1][30][1] ,
         \s_mux1_signals[1][30][0] , \s_mux1_signals[2][0][31] ,
         \s_mux1_signals[2][0][30] , \s_mux1_signals[2][0][29] ,
         \s_mux1_signals[2][0][28] , \s_mux1_signals[2][0][27] ,
         \s_mux1_signals[2][0][26] , \s_mux1_signals[2][0][25] ,
         \s_mux1_signals[2][0][24] , \s_mux1_signals[2][0][23] ,
         \s_mux1_signals[2][0][22] , \s_mux1_signals[2][0][21] ,
         \s_mux1_signals[2][0][20] , \s_mux1_signals[2][0][19] ,
         \s_mux1_signals[2][0][18] , \s_mux1_signals[2][0][17] ,
         \s_mux1_signals[2][0][16] , \s_mux1_signals[2][0][15] ,
         \s_mux1_signals[2][0][14] , \s_mux1_signals[2][0][13] ,
         \s_mux1_signals[2][0][12] , \s_mux1_signals[2][0][11] ,
         \s_mux1_signals[2][0][10] , \s_mux1_signals[2][0][9] ,
         \s_mux1_signals[2][0][8] , \s_mux1_signals[2][0][7] ,
         \s_mux1_signals[2][0][6] , \s_mux1_signals[2][0][5] ,
         \s_mux1_signals[2][0][4] , \s_mux1_signals[2][0][3] ,
         \s_mux1_signals[2][0][2] , \s_mux1_signals[2][0][1] ,
         \s_mux1_signals[2][0][0] , \s_mux1_signals[2][4][31] ,
         \s_mux1_signals[2][4][30] , \s_mux1_signals[2][4][29] ,
         \s_mux1_signals[2][4][28] , \s_mux1_signals[2][4][27] ,
         \s_mux1_signals[2][4][26] , \s_mux1_signals[2][4][25] ,
         \s_mux1_signals[2][4][24] , \s_mux1_signals[2][4][23] ,
         \s_mux1_signals[2][4][22] , \s_mux1_signals[2][4][21] ,
         \s_mux1_signals[2][4][20] , \s_mux1_signals[2][4][19] ,
         \s_mux1_signals[2][4][18] , \s_mux1_signals[2][4][17] ,
         \s_mux1_signals[2][4][16] , \s_mux1_signals[2][4][15] ,
         \s_mux1_signals[2][4][14] , \s_mux1_signals[2][4][13] ,
         \s_mux1_signals[2][4][12] , \s_mux1_signals[2][4][11] ,
         \s_mux1_signals[2][4][10] , \s_mux1_signals[2][4][9] ,
         \s_mux1_signals[2][4][8] , \s_mux1_signals[2][4][7] ,
         \s_mux1_signals[2][4][6] , \s_mux1_signals[2][4][5] ,
         \s_mux1_signals[2][4][4] , \s_mux1_signals[2][4][3] ,
         \s_mux1_signals[2][4][2] , \s_mux1_signals[2][4][1] ,
         \s_mux1_signals[2][4][0] , \s_mux1_signals[2][8][31] ,
         \s_mux1_signals[2][8][30] , \s_mux1_signals[2][8][29] ,
         \s_mux1_signals[2][8][28] , \s_mux1_signals[2][8][27] ,
         \s_mux1_signals[2][8][26] , \s_mux1_signals[2][8][25] ,
         \s_mux1_signals[2][8][24] , \s_mux1_signals[2][8][23] ,
         \s_mux1_signals[2][8][22] , \s_mux1_signals[2][8][21] ,
         \s_mux1_signals[2][8][20] , \s_mux1_signals[2][8][19] ,
         \s_mux1_signals[2][8][18] , \s_mux1_signals[2][8][17] ,
         \s_mux1_signals[2][8][16] , \s_mux1_signals[2][8][15] ,
         \s_mux1_signals[2][8][14] , \s_mux1_signals[2][8][13] ,
         \s_mux1_signals[2][8][12] , \s_mux1_signals[2][8][11] ,
         \s_mux1_signals[2][8][10] , \s_mux1_signals[2][8][9] ,
         \s_mux1_signals[2][8][8] , \s_mux1_signals[2][8][7] ,
         \s_mux1_signals[2][8][6] , \s_mux1_signals[2][8][5] ,
         \s_mux1_signals[2][8][4] , \s_mux1_signals[2][8][3] ,
         \s_mux1_signals[2][8][2] , \s_mux1_signals[2][8][1] ,
         \s_mux1_signals[2][8][0] , \s_mux1_signals[2][12][31] ,
         \s_mux1_signals[2][12][30] , \s_mux1_signals[2][12][29] ,
         \s_mux1_signals[2][12][28] , \s_mux1_signals[2][12][27] ,
         \s_mux1_signals[2][12][26] , \s_mux1_signals[2][12][25] ,
         \s_mux1_signals[2][12][24] , \s_mux1_signals[2][12][23] ,
         \s_mux1_signals[2][12][22] , \s_mux1_signals[2][12][21] ,
         \s_mux1_signals[2][12][20] , \s_mux1_signals[2][12][19] ,
         \s_mux1_signals[2][12][18] , \s_mux1_signals[2][12][17] ,
         \s_mux1_signals[2][12][16] , \s_mux1_signals[2][12][15] ,
         \s_mux1_signals[2][12][14] , \s_mux1_signals[2][12][13] ,
         \s_mux1_signals[2][12][12] , \s_mux1_signals[2][12][11] ,
         \s_mux1_signals[2][12][10] , \s_mux1_signals[2][12][9] ,
         \s_mux1_signals[2][12][8] , \s_mux1_signals[2][12][7] ,
         \s_mux1_signals[2][12][6] , \s_mux1_signals[2][12][5] ,
         \s_mux1_signals[2][12][4] , \s_mux1_signals[2][12][3] ,
         \s_mux1_signals[2][12][2] , \s_mux1_signals[2][12][1] ,
         \s_mux1_signals[2][12][0] , \s_mux1_signals[2][16][31] ,
         \s_mux1_signals[2][16][30] , \s_mux1_signals[2][16][29] ,
         \s_mux1_signals[2][16][28] , \s_mux1_signals[2][16][27] ,
         \s_mux1_signals[2][16][26] , \s_mux1_signals[2][16][25] ,
         \s_mux1_signals[2][16][24] , \s_mux1_signals[2][16][23] ,
         \s_mux1_signals[2][16][22] , \s_mux1_signals[2][16][21] ,
         \s_mux1_signals[2][16][20] , \s_mux1_signals[2][16][19] ,
         \s_mux1_signals[2][16][18] , \s_mux1_signals[2][16][17] ,
         \s_mux1_signals[2][16][16] , \s_mux1_signals[2][16][15] ,
         \s_mux1_signals[2][16][14] , \s_mux1_signals[2][16][13] ,
         \s_mux1_signals[2][16][12] , \s_mux1_signals[2][16][11] ,
         \s_mux1_signals[2][16][10] , \s_mux1_signals[2][16][9] ,
         \s_mux1_signals[2][16][8] , \s_mux1_signals[2][16][7] ,
         \s_mux1_signals[2][16][6] , \s_mux1_signals[2][16][5] ,
         \s_mux1_signals[2][16][4] , \s_mux1_signals[2][16][3] ,
         \s_mux1_signals[2][16][2] , \s_mux1_signals[2][16][1] ,
         \s_mux1_signals[2][16][0] , \s_mux1_signals[2][20][31] ,
         \s_mux1_signals[2][20][30] , \s_mux1_signals[2][20][29] ,
         \s_mux1_signals[2][20][28] , \s_mux1_signals[2][20][27] ,
         \s_mux1_signals[2][20][26] , \s_mux1_signals[2][20][25] ,
         \s_mux1_signals[2][20][24] , \s_mux1_signals[2][20][23] ,
         \s_mux1_signals[2][20][22] , \s_mux1_signals[2][20][21] ,
         \s_mux1_signals[2][20][20] , \s_mux1_signals[2][20][19] ,
         \s_mux1_signals[2][20][18] , \s_mux1_signals[2][20][17] ,
         \s_mux1_signals[2][20][16] , \s_mux1_signals[2][20][15] ,
         \s_mux1_signals[2][20][14] , \s_mux1_signals[2][20][13] ,
         \s_mux1_signals[2][20][12] , \s_mux1_signals[2][20][11] ,
         \s_mux1_signals[2][20][10] , \s_mux1_signals[2][20][9] ,
         \s_mux1_signals[2][20][8] , \s_mux1_signals[2][20][7] ,
         \s_mux1_signals[2][20][6] , \s_mux1_signals[2][20][5] ,
         \s_mux1_signals[2][20][4] , \s_mux1_signals[2][20][3] ,
         \s_mux1_signals[2][20][2] , \s_mux1_signals[2][20][1] ,
         \s_mux1_signals[2][20][0] , \s_mux1_signals[2][24][31] ,
         \s_mux1_signals[2][24][30] , \s_mux1_signals[2][24][29] ,
         \s_mux1_signals[2][24][28] , \s_mux1_signals[2][24][27] ,
         \s_mux1_signals[2][24][26] , \s_mux1_signals[2][24][25] ,
         \s_mux1_signals[2][24][24] , \s_mux1_signals[2][24][23] ,
         \s_mux1_signals[2][24][22] , \s_mux1_signals[2][24][21] ,
         \s_mux1_signals[2][24][20] , \s_mux1_signals[2][24][19] ,
         \s_mux1_signals[2][24][18] , \s_mux1_signals[2][24][17] ,
         \s_mux1_signals[2][24][16] , \s_mux1_signals[2][24][15] ,
         \s_mux1_signals[2][24][14] , \s_mux1_signals[2][24][13] ,
         \s_mux1_signals[2][24][12] , \s_mux1_signals[2][24][11] ,
         \s_mux1_signals[2][24][10] , \s_mux1_signals[2][24][9] ,
         \s_mux1_signals[2][24][8] , \s_mux1_signals[2][24][7] ,
         \s_mux1_signals[2][24][6] , \s_mux1_signals[2][24][5] ,
         \s_mux1_signals[2][24][4] , \s_mux1_signals[2][24][3] ,
         \s_mux1_signals[2][24][2] , \s_mux1_signals[2][24][1] ,
         \s_mux1_signals[2][24][0] , \s_mux1_signals[2][28][31] ,
         \s_mux1_signals[2][28][30] , \s_mux1_signals[2][28][29] ,
         \s_mux1_signals[2][28][28] , \s_mux1_signals[2][28][27] ,
         \s_mux1_signals[2][28][26] , \s_mux1_signals[2][28][25] ,
         \s_mux1_signals[2][28][24] , \s_mux1_signals[2][28][23] ,
         \s_mux1_signals[2][28][22] , \s_mux1_signals[2][28][21] ,
         \s_mux1_signals[2][28][20] , \s_mux1_signals[2][28][19] ,
         \s_mux1_signals[2][28][18] , \s_mux1_signals[2][28][17] ,
         \s_mux1_signals[2][28][16] , \s_mux1_signals[2][28][15] ,
         \s_mux1_signals[2][28][14] , \s_mux1_signals[2][28][13] ,
         \s_mux1_signals[2][28][12] , \s_mux1_signals[2][28][11] ,
         \s_mux1_signals[2][28][10] , \s_mux1_signals[2][28][9] ,
         \s_mux1_signals[2][28][8] , \s_mux1_signals[2][28][7] ,
         \s_mux1_signals[2][28][6] , \s_mux1_signals[2][28][5] ,
         \s_mux1_signals[2][28][4] , \s_mux1_signals[2][28][3] ,
         \s_mux1_signals[2][28][2] , \s_mux1_signals[2][28][1] ,
         \s_mux1_signals[2][28][0] , \s_mux1_signals[3][0][31] ,
         \s_mux1_signals[3][0][30] , \s_mux1_signals[3][0][29] ,
         \s_mux1_signals[3][0][28] , \s_mux1_signals[3][0][27] ,
         \s_mux1_signals[3][0][26] , \s_mux1_signals[3][0][25] ,
         \s_mux1_signals[3][0][24] , \s_mux1_signals[3][0][23] ,
         \s_mux1_signals[3][0][22] , \s_mux1_signals[3][0][21] ,
         \s_mux1_signals[3][0][20] , \s_mux1_signals[3][0][19] ,
         \s_mux1_signals[3][0][18] , \s_mux1_signals[3][0][17] ,
         \s_mux1_signals[3][0][16] , \s_mux1_signals[3][0][15] ,
         \s_mux1_signals[3][0][14] , \s_mux1_signals[3][0][13] ,
         \s_mux1_signals[3][0][12] , \s_mux1_signals[3][0][11] ,
         \s_mux1_signals[3][0][10] , \s_mux1_signals[3][0][9] ,
         \s_mux1_signals[3][0][8] , \s_mux1_signals[3][0][7] ,
         \s_mux1_signals[3][0][6] , \s_mux1_signals[3][0][5] ,
         \s_mux1_signals[3][0][4] , \s_mux1_signals[3][0][3] ,
         \s_mux1_signals[3][0][2] , \s_mux1_signals[3][0][1] ,
         \s_mux1_signals[3][0][0] , \s_mux1_signals[3][8][31] ,
         \s_mux1_signals[3][8][30] , \s_mux1_signals[3][8][29] ,
         \s_mux1_signals[3][8][28] , \s_mux1_signals[3][8][27] ,
         \s_mux1_signals[3][8][26] , \s_mux1_signals[3][8][25] ,
         \s_mux1_signals[3][8][24] , \s_mux1_signals[3][8][23] ,
         \s_mux1_signals[3][8][22] , \s_mux1_signals[3][8][21] ,
         \s_mux1_signals[3][8][20] , \s_mux1_signals[3][8][19] ,
         \s_mux1_signals[3][8][18] , \s_mux1_signals[3][8][17] ,
         \s_mux1_signals[3][8][16] , \s_mux1_signals[3][8][15] ,
         \s_mux1_signals[3][8][14] , \s_mux1_signals[3][8][13] ,
         \s_mux1_signals[3][8][12] , \s_mux1_signals[3][8][11] ,
         \s_mux1_signals[3][8][10] , \s_mux1_signals[3][8][9] ,
         \s_mux1_signals[3][8][8] , \s_mux1_signals[3][8][7] ,
         \s_mux1_signals[3][8][6] , \s_mux1_signals[3][8][5] ,
         \s_mux1_signals[3][8][4] , \s_mux1_signals[3][8][3] ,
         \s_mux1_signals[3][8][2] , \s_mux1_signals[3][8][1] ,
         \s_mux1_signals[3][8][0] , \s_mux1_signals[3][16][31] ,
         \s_mux1_signals[3][16][30] , \s_mux1_signals[3][16][29] ,
         \s_mux1_signals[3][16][28] , \s_mux1_signals[3][16][27] ,
         \s_mux1_signals[3][16][26] , \s_mux1_signals[3][16][25] ,
         \s_mux1_signals[3][16][24] , \s_mux1_signals[3][16][23] ,
         \s_mux1_signals[3][16][22] , \s_mux1_signals[3][16][21] ,
         \s_mux1_signals[3][16][20] , \s_mux1_signals[3][16][19] ,
         \s_mux1_signals[3][16][18] , \s_mux1_signals[3][16][17] ,
         \s_mux1_signals[3][16][16] , \s_mux1_signals[3][16][15] ,
         \s_mux1_signals[3][16][14] , \s_mux1_signals[3][16][13] ,
         \s_mux1_signals[3][16][12] , \s_mux1_signals[3][16][11] ,
         \s_mux1_signals[3][16][10] , \s_mux1_signals[3][16][9] ,
         \s_mux1_signals[3][16][8] , \s_mux1_signals[3][16][7] ,
         \s_mux1_signals[3][16][6] , \s_mux1_signals[3][16][5] ,
         \s_mux1_signals[3][16][4] , \s_mux1_signals[3][16][3] ,
         \s_mux1_signals[3][16][2] , \s_mux1_signals[3][16][1] ,
         \s_mux1_signals[3][16][0] , \s_mux1_signals[3][24][31] ,
         \s_mux1_signals[3][24][30] , \s_mux1_signals[3][24][29] ,
         \s_mux1_signals[3][24][28] , \s_mux1_signals[3][24][27] ,
         \s_mux1_signals[3][24][26] , \s_mux1_signals[3][24][25] ,
         \s_mux1_signals[3][24][24] , \s_mux1_signals[3][24][23] ,
         \s_mux1_signals[3][24][22] , \s_mux1_signals[3][24][21] ,
         \s_mux1_signals[3][24][20] , \s_mux1_signals[3][24][19] ,
         \s_mux1_signals[3][24][18] , \s_mux1_signals[3][24][17] ,
         \s_mux1_signals[3][24][16] , \s_mux1_signals[3][24][15] ,
         \s_mux1_signals[3][24][14] , \s_mux1_signals[3][24][13] ,
         \s_mux1_signals[3][24][12] , \s_mux1_signals[3][24][11] ,
         \s_mux1_signals[3][24][10] , \s_mux1_signals[3][24][9] ,
         \s_mux1_signals[3][24][8] , \s_mux1_signals[3][24][7] ,
         \s_mux1_signals[3][24][6] , \s_mux1_signals[3][24][5] ,
         \s_mux1_signals[3][24][4] , \s_mux1_signals[3][24][3] ,
         \s_mux1_signals[3][24][2] , \s_mux1_signals[3][24][1] ,
         \s_mux1_signals[3][24][0] , \s_mux1_signals[4][0][31] ,
         \s_mux1_signals[4][0][30] , \s_mux1_signals[4][0][29] ,
         \s_mux1_signals[4][0][28] , \s_mux1_signals[4][0][27] ,
         \s_mux1_signals[4][0][26] , \s_mux1_signals[4][0][25] ,
         \s_mux1_signals[4][0][24] , \s_mux1_signals[4][0][23] ,
         \s_mux1_signals[4][0][22] , \s_mux1_signals[4][0][21] ,
         \s_mux1_signals[4][0][20] , \s_mux1_signals[4][0][19] ,
         \s_mux1_signals[4][0][18] , \s_mux1_signals[4][0][17] ,
         \s_mux1_signals[4][0][16] , \s_mux1_signals[4][0][15] ,
         \s_mux1_signals[4][0][14] , \s_mux1_signals[4][0][13] ,
         \s_mux1_signals[4][0][12] , \s_mux1_signals[4][0][11] ,
         \s_mux1_signals[4][0][10] , \s_mux1_signals[4][0][9] ,
         \s_mux1_signals[4][0][8] , \s_mux1_signals[4][0][7] ,
         \s_mux1_signals[4][0][6] , \s_mux1_signals[4][0][5] ,
         \s_mux1_signals[4][0][4] , \s_mux1_signals[4][0][3] ,
         \s_mux1_signals[4][0][2] , \s_mux1_signals[4][0][1] ,
         \s_mux1_signals[4][0][0] , \s_mux1_signals[4][16][31] ,
         \s_mux1_signals[4][16][30] , \s_mux1_signals[4][16][29] ,
         \s_mux1_signals[4][16][28] , \s_mux1_signals[4][16][27] ,
         \s_mux1_signals[4][16][26] , \s_mux1_signals[4][16][25] ,
         \s_mux1_signals[4][16][24] , \s_mux1_signals[4][16][23] ,
         \s_mux1_signals[4][16][22] , \s_mux1_signals[4][16][21] ,
         \s_mux1_signals[4][16][20] , \s_mux1_signals[4][16][19] ,
         \s_mux1_signals[4][16][18] , \s_mux1_signals[4][16][17] ,
         \s_mux1_signals[4][16][16] , \s_mux1_signals[4][16][15] ,
         \s_mux1_signals[4][16][14] , \s_mux1_signals[4][16][13] ,
         \s_mux1_signals[4][16][12] , \s_mux1_signals[4][16][11] ,
         \s_mux1_signals[4][16][10] , \s_mux1_signals[4][16][9] ,
         \s_mux1_signals[4][16][8] , \s_mux1_signals[4][16][7] ,
         \s_mux1_signals[4][16][6] , \s_mux1_signals[4][16][5] ,
         \s_mux1_signals[4][16][4] , \s_mux1_signals[4][16][3] ,
         \s_mux1_signals[4][16][2] , \s_mux1_signals[4][16][1] ,
         \s_mux1_signals[4][16][0] , n2, n4, n9, n21, n22, n23, n24, n25, n26,
         n27, n28, n29, n30, n31, n32, n33, n34, n35, n36, n37, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68,
         n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82,
         n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n97, n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108,
         n109, n110, n111, n112, n113, n114, n115, n116, n117, n118, n119;
  wire   [31:1] s_load_Fdec_Tregs;
  wire   [4:0] s_addrRd1_Fei_Tmux;
  wire   [4:0] s_addrRd2_Fei_Tmux;
  wire   SYNOPSYS_UNCONNECTED__0;

  INV_X2 U5 ( .A(RF_clk), .ZN(n9) );
  Decoder_DEC_NBIT5 WR_DEC ( .DEC_address(RF_AddrWr), .DEC_enable(s_wr_enable), 
        .DEC_output({s_load_Fdec_Tregs, SYNOPSYS_UNCONNECTED__0}) );
  Enable_Interface_NBIT_DATA5_0 RD1_EI ( .EI_datain(RF_AddrRd1), .EI_enable(
        s_rd1_enable), .EI_dataout({s_addrRd1_Fei_Tmux[4:1], n4}) );
  Enable_Interface_NBIT_DATA5_1 RD2_EI ( .EI_datain(RF_AddrRd2), .EI_enable(
        s_rd2_enable), .EI_dataout({s_addrRd2_Fei_Tmux[4:1], n2}) );
  NRegister_N32_32 R0_0 ( .clk(n9), .reset(n119), .data_in({1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .enable(n116), .load(1'b0), .data_out(
        {\s_mux2_signals[0][0][31] , \s_mux2_signals[0][0][30] , 
        \s_mux2_signals[0][0][29] , \s_mux2_signals[0][0][28] , 
        \s_mux2_signals[0][0][27] , \s_mux2_signals[0][0][26] , 
        \s_mux2_signals[0][0][25] , \s_mux2_signals[0][0][24] , 
        \s_mux2_signals[0][0][23] , \s_mux2_signals[0][0][22] , 
        \s_mux2_signals[0][0][21] , \s_mux2_signals[0][0][20] , 
        \s_mux2_signals[0][0][19] , \s_mux2_signals[0][0][18] , 
        \s_mux2_signals[0][0][17] , \s_mux2_signals[0][0][16] , 
        \s_mux2_signals[0][0][15] , \s_mux2_signals[0][0][14] , 
        \s_mux2_signals[0][0][13] , \s_mux2_signals[0][0][12] , 
        \s_mux2_signals[0][0][11] , \s_mux2_signals[0][0][10] , 
        \s_mux2_signals[0][0][9] , \s_mux2_signals[0][0][8] , 
        \s_mux2_signals[0][0][7] , \s_mux2_signals[0][0][6] , 
        \s_mux2_signals[0][0][5] , \s_mux2_signals[0][0][4] , 
        \s_mux2_signals[0][0][3] , \s_mux2_signals[0][0][2] , 
        \s_mux2_signals[0][0][1] , \s_mux2_signals[0][0][0] }) );
  NRegister_N32_31 Ri_1 ( .clk(n9), .reset(n119), .data_in({RF_data_in[31], 
        n112, n111, n110, n109, n108, n107, n104, n101, n98, n97, n94, n91, 
        n88, n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, 
        n46, n43, n40, n37, n36}), .enable(n116), .load(s_load_Fdec_Tregs[1]), 
        .data_out({\s_mux2_signals[0][1][31] , \s_mux2_signals[0][1][30] , 
        \s_mux2_signals[0][1][29] , \s_mux2_signals[0][1][28] , 
        \s_mux2_signals[0][1][27] , \s_mux2_signals[0][1][26] , 
        \s_mux2_signals[0][1][25] , \s_mux2_signals[0][1][24] , 
        \s_mux2_signals[0][1][23] , \s_mux2_signals[0][1][22] , 
        \s_mux2_signals[0][1][21] , \s_mux2_signals[0][1][20] , 
        \s_mux2_signals[0][1][19] , \s_mux2_signals[0][1][18] , 
        \s_mux2_signals[0][1][17] , \s_mux2_signals[0][1][16] , 
        \s_mux2_signals[0][1][15] , \s_mux2_signals[0][1][14] , 
        \s_mux2_signals[0][1][13] , \s_mux2_signals[0][1][12] , 
        \s_mux2_signals[0][1][11] , \s_mux2_signals[0][1][10] , 
        \s_mux2_signals[0][1][9] , \s_mux2_signals[0][1][8] , 
        \s_mux2_signals[0][1][7] , \s_mux2_signals[0][1][6] , 
        \s_mux2_signals[0][1][5] , \s_mux2_signals[0][1][4] , 
        \s_mux2_signals[0][1][3] , \s_mux2_signals[0][1][2] , 
        \s_mux2_signals[0][1][1] , \s_mux2_signals[0][1][0] }) );
  NRegister_N32_30 Ri_2 ( .clk(n9), .reset(n117), .data_in({n113, 
        RF_data_in[30:26], n105, n102, n99, RF_data_in[22], n95, n92, n89, n86, 
        n83, n80, n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, n44, 
        n41, n38, RF_data_in[1:0]}), .enable(n114), .load(s_load_Fdec_Tregs[2]), .data_out({\s_mux2_signals[0][2][31] , \s_mux2_signals[0][2][30] , 
        \s_mux2_signals[0][2][29] , \s_mux2_signals[0][2][28] , 
        \s_mux2_signals[0][2][27] , \s_mux2_signals[0][2][26] , 
        \s_mux2_signals[0][2][25] , \s_mux2_signals[0][2][24] , 
        \s_mux2_signals[0][2][23] , \s_mux2_signals[0][2][22] , 
        \s_mux2_signals[0][2][21] , \s_mux2_signals[0][2][20] , 
        \s_mux2_signals[0][2][19] , \s_mux2_signals[0][2][18] , 
        \s_mux2_signals[0][2][17] , \s_mux2_signals[0][2][16] , 
        \s_mux2_signals[0][2][15] , \s_mux2_signals[0][2][14] , 
        \s_mux2_signals[0][2][13] , \s_mux2_signals[0][2][12] , 
        \s_mux2_signals[0][2][11] , \s_mux2_signals[0][2][10] , 
        \s_mux2_signals[0][2][9] , \s_mux2_signals[0][2][8] , 
        \s_mux2_signals[0][2][7] , \s_mux2_signals[0][2][6] , 
        \s_mux2_signals[0][2][5] , \s_mux2_signals[0][2][4] , 
        \s_mux2_signals[0][2][3] , \s_mux2_signals[0][2][2] , 
        \s_mux2_signals[0][2][1] , \s_mux2_signals[0][2][0] }) );
  NRegister_N32_29 Ri_3 ( .clk(n9), .reset(n117), .data_in({n113, n112, n111, 
        n110, n109, n108, n105, n102, n99, n98, n95, n92, n89, n86, n83, n80, 
        n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, n44, n41, n38, 
        n37, n36}), .enable(n114), .load(s_load_Fdec_Tregs[3]), .data_out({
        \s_mux2_signals[0][3][31] , \s_mux2_signals[0][3][30] , 
        \s_mux2_signals[0][3][29] , \s_mux2_signals[0][3][28] , 
        \s_mux2_signals[0][3][27] , \s_mux2_signals[0][3][26] , 
        \s_mux2_signals[0][3][25] , \s_mux2_signals[0][3][24] , 
        \s_mux2_signals[0][3][23] , \s_mux2_signals[0][3][22] , 
        \s_mux2_signals[0][3][21] , \s_mux2_signals[0][3][20] , 
        \s_mux2_signals[0][3][19] , \s_mux2_signals[0][3][18] , 
        \s_mux2_signals[0][3][17] , \s_mux2_signals[0][3][16] , 
        \s_mux2_signals[0][3][15] , \s_mux2_signals[0][3][14] , 
        \s_mux2_signals[0][3][13] , \s_mux2_signals[0][3][12] , 
        \s_mux2_signals[0][3][11] , \s_mux2_signals[0][3][10] , 
        \s_mux2_signals[0][3][9] , \s_mux2_signals[0][3][8] , 
        \s_mux2_signals[0][3][7] , \s_mux2_signals[0][3][6] , 
        \s_mux2_signals[0][3][5] , \s_mux2_signals[0][3][4] , 
        \s_mux2_signals[0][3][3] , \s_mux2_signals[0][3][2] , 
        \s_mux2_signals[0][3][1] , \s_mux2_signals[0][3][0] }) );
  NRegister_N32_28 Ri_4 ( .clk(n9), .reset(n117), .data_in({n113, n112, n111, 
        n110, n109, n108, n105, n102, n99, n98, n95, n92, n89, n86, n83, n80, 
        n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, n44, n41, n38, 
        n37, n36}), .enable(n114), .load(s_load_Fdec_Tregs[4]), .data_out({
        \s_mux2_signals[0][4][31] , \s_mux2_signals[0][4][30] , 
        \s_mux2_signals[0][4][29] , \s_mux2_signals[0][4][28] , 
        \s_mux2_signals[0][4][27] , \s_mux2_signals[0][4][26] , 
        \s_mux2_signals[0][4][25] , \s_mux2_signals[0][4][24] , 
        \s_mux2_signals[0][4][23] , \s_mux2_signals[0][4][22] , 
        \s_mux2_signals[0][4][21] , \s_mux2_signals[0][4][20] , 
        \s_mux2_signals[0][4][19] , \s_mux2_signals[0][4][18] , 
        \s_mux2_signals[0][4][17] , \s_mux2_signals[0][4][16] , 
        \s_mux2_signals[0][4][15] , \s_mux2_signals[0][4][14] , 
        \s_mux2_signals[0][4][13] , \s_mux2_signals[0][4][12] , 
        \s_mux2_signals[0][4][11] , \s_mux2_signals[0][4][10] , 
        \s_mux2_signals[0][4][9] , \s_mux2_signals[0][4][8] , 
        \s_mux2_signals[0][4][7] , \s_mux2_signals[0][4][6] , 
        \s_mux2_signals[0][4][5] , \s_mux2_signals[0][4][4] , 
        \s_mux2_signals[0][4][3] , \s_mux2_signals[0][4][2] , 
        \s_mux2_signals[0][4][1] , \s_mux2_signals[0][4][0] }) );
  NRegister_N32_27 Ri_5 ( .clk(n9), .reset(n117), .data_in({n113, n112, n111, 
        n110, n109, n108, n105, n102, n99, n98, n95, n92, n89, n86, n83, n80, 
        n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, n44, n41, n38, 
        n37, n36}), .enable(n114), .load(s_load_Fdec_Tregs[5]), .data_out({
        \s_mux2_signals[0][5][31] , \s_mux2_signals[0][5][30] , 
        \s_mux2_signals[0][5][29] , \s_mux2_signals[0][5][28] , 
        \s_mux2_signals[0][5][27] , \s_mux2_signals[0][5][26] , 
        \s_mux2_signals[0][5][25] , \s_mux2_signals[0][5][24] , 
        \s_mux2_signals[0][5][23] , \s_mux2_signals[0][5][22] , 
        \s_mux2_signals[0][5][21] , \s_mux2_signals[0][5][20] , 
        \s_mux2_signals[0][5][19] , \s_mux2_signals[0][5][18] , 
        \s_mux2_signals[0][5][17] , \s_mux2_signals[0][5][16] , 
        \s_mux2_signals[0][5][15] , \s_mux2_signals[0][5][14] , 
        \s_mux2_signals[0][5][13] , \s_mux2_signals[0][5][12] , 
        \s_mux2_signals[0][5][11] , \s_mux2_signals[0][5][10] , 
        \s_mux2_signals[0][5][9] , \s_mux2_signals[0][5][8] , 
        \s_mux2_signals[0][5][7] , \s_mux2_signals[0][5][6] , 
        \s_mux2_signals[0][5][5] , \s_mux2_signals[0][5][4] , 
        \s_mux2_signals[0][5][3] , \s_mux2_signals[0][5][2] , 
        \s_mux2_signals[0][5][1] , \s_mux2_signals[0][5][0] }) );
  NRegister_N32_26 Ri_6 ( .clk(n9), .reset(n117), .data_in({n113, n112, n111, 
        n110, n109, n108, n105, n102, n99, n98, n95, n92, n89, n86, n83, n80, 
        n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, n44, n41, n38, 
        n37, n36}), .enable(n114), .load(s_load_Fdec_Tregs[6]), .data_out({
        \s_mux2_signals[0][6][31] , \s_mux2_signals[0][6][30] , 
        \s_mux2_signals[0][6][29] , \s_mux2_signals[0][6][28] , 
        \s_mux2_signals[0][6][27] , \s_mux2_signals[0][6][26] , 
        \s_mux2_signals[0][6][25] , \s_mux2_signals[0][6][24] , 
        \s_mux2_signals[0][6][23] , \s_mux2_signals[0][6][22] , 
        \s_mux2_signals[0][6][21] , \s_mux2_signals[0][6][20] , 
        \s_mux2_signals[0][6][19] , \s_mux2_signals[0][6][18] , 
        \s_mux2_signals[0][6][17] , \s_mux2_signals[0][6][16] , 
        \s_mux2_signals[0][6][15] , \s_mux2_signals[0][6][14] , 
        \s_mux2_signals[0][6][13] , \s_mux2_signals[0][6][12] , 
        \s_mux2_signals[0][6][11] , \s_mux2_signals[0][6][10] , 
        \s_mux2_signals[0][6][9] , \s_mux2_signals[0][6][8] , 
        \s_mux2_signals[0][6][7] , \s_mux2_signals[0][6][6] , 
        \s_mux2_signals[0][6][5] , \s_mux2_signals[0][6][4] , 
        \s_mux2_signals[0][6][3] , \s_mux2_signals[0][6][2] , 
        \s_mux2_signals[0][6][1] , \s_mux2_signals[0][6][0] }) );
  NRegister_N32_25 Ri_7 ( .clk(n9), .reset(n117), .data_in({n113, n112, n111, 
        n110, n109, n108, n105, n102, n99, n98, n95, n92, n89, n86, n83, n80, 
        n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, n44, n41, n38, 
        n37, n36}), .enable(n114), .load(s_load_Fdec_Tregs[7]), .data_out({
        \s_mux2_signals[0][7][31] , \s_mux2_signals[0][7][30] , 
        \s_mux2_signals[0][7][29] , \s_mux2_signals[0][7][28] , 
        \s_mux2_signals[0][7][27] , \s_mux2_signals[0][7][26] , 
        \s_mux2_signals[0][7][25] , \s_mux2_signals[0][7][24] , 
        \s_mux2_signals[0][7][23] , \s_mux2_signals[0][7][22] , 
        \s_mux2_signals[0][7][21] , \s_mux2_signals[0][7][20] , 
        \s_mux2_signals[0][7][19] , \s_mux2_signals[0][7][18] , 
        \s_mux2_signals[0][7][17] , \s_mux2_signals[0][7][16] , 
        \s_mux2_signals[0][7][15] , \s_mux2_signals[0][7][14] , 
        \s_mux2_signals[0][7][13] , \s_mux2_signals[0][7][12] , 
        \s_mux2_signals[0][7][11] , \s_mux2_signals[0][7][10] , 
        \s_mux2_signals[0][7][9] , \s_mux2_signals[0][7][8] , 
        \s_mux2_signals[0][7][7] , \s_mux2_signals[0][7][6] , 
        \s_mux2_signals[0][7][5] , \s_mux2_signals[0][7][4] , 
        \s_mux2_signals[0][7][3] , \s_mux2_signals[0][7][2] , 
        \s_mux2_signals[0][7][1] , \s_mux2_signals[0][7][0] }) );
  NRegister_N32_24 Ri_8 ( .clk(n9), .reset(n119), .data_in({RF_data_in[31], 
        n112, n111, n110, n109, n108, n107, n104, n101, n98, n97, n94, n91, 
        n88, n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, 
        n46, n43, n40, n37, n36}), .enable(n116), .load(s_load_Fdec_Tregs[8]), 
        .data_out({\s_mux2_signals[0][8][31] , \s_mux2_signals[0][8][30] , 
        \s_mux2_signals[0][8][29] , \s_mux2_signals[0][8][28] , 
        \s_mux2_signals[0][8][27] , \s_mux2_signals[0][8][26] , 
        \s_mux2_signals[0][8][25] , \s_mux2_signals[0][8][24] , 
        \s_mux2_signals[0][8][23] , \s_mux2_signals[0][8][22] , 
        \s_mux2_signals[0][8][21] , \s_mux2_signals[0][8][20] , 
        \s_mux2_signals[0][8][19] , \s_mux2_signals[0][8][18] , 
        \s_mux2_signals[0][8][17] , \s_mux2_signals[0][8][16] , 
        \s_mux2_signals[0][8][15] , \s_mux2_signals[0][8][14] , 
        \s_mux2_signals[0][8][13] , \s_mux2_signals[0][8][12] , 
        \s_mux2_signals[0][8][11] , \s_mux2_signals[0][8][10] , 
        \s_mux2_signals[0][8][9] , \s_mux2_signals[0][8][8] , 
        \s_mux2_signals[0][8][7] , \s_mux2_signals[0][8][6] , 
        \s_mux2_signals[0][8][5] , \s_mux2_signals[0][8][4] , 
        \s_mux2_signals[0][8][3] , \s_mux2_signals[0][8][2] , 
        \s_mux2_signals[0][8][1] , \s_mux2_signals[0][8][0] }) );
  NRegister_N32_23 Ri_9 ( .clk(n9), .reset(n117), .data_in({n113, 
        RF_data_in[30:26], n105, n102, n99, RF_data_in[22], n95, n92, n89, n86, 
        n83, n80, n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, n44, 
        n41, n38, RF_data_in[1:0]}), .enable(n114), .load(s_load_Fdec_Tregs[9]), .data_out({\s_mux2_signals[0][9][31] , \s_mux2_signals[0][9][30] , 
        \s_mux2_signals[0][9][29] , \s_mux2_signals[0][9][28] , 
        \s_mux2_signals[0][9][27] , \s_mux2_signals[0][9][26] , 
        \s_mux2_signals[0][9][25] , \s_mux2_signals[0][9][24] , 
        \s_mux2_signals[0][9][23] , \s_mux2_signals[0][9][22] , 
        \s_mux2_signals[0][9][21] , \s_mux2_signals[0][9][20] , 
        \s_mux2_signals[0][9][19] , \s_mux2_signals[0][9][18] , 
        \s_mux2_signals[0][9][17] , \s_mux2_signals[0][9][16] , 
        \s_mux2_signals[0][9][15] , \s_mux2_signals[0][9][14] , 
        \s_mux2_signals[0][9][13] , \s_mux2_signals[0][9][12] , 
        \s_mux2_signals[0][9][11] , \s_mux2_signals[0][9][10] , 
        \s_mux2_signals[0][9][9] , \s_mux2_signals[0][9][8] , 
        \s_mux2_signals[0][9][7] , \s_mux2_signals[0][9][6] , 
        \s_mux2_signals[0][9][5] , \s_mux2_signals[0][9][4] , 
        \s_mux2_signals[0][9][3] , \s_mux2_signals[0][9][2] , 
        \s_mux2_signals[0][9][1] , \s_mux2_signals[0][9][0] }) );
  NRegister_N32_22 Ri_10 ( .clk(n9), .reset(n117), .data_in({n113, 
        RF_data_in[30:26], n105, n102, n99, RF_data_in[22], n95, n92, n89, n86, 
        n83, n80, n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, n44, 
        n41, n38, RF_data_in[1:0]}), .enable(n114), .load(
        s_load_Fdec_Tregs[10]), .data_out({\s_mux2_signals[0][10][31] , 
        \s_mux2_signals[0][10][30] , \s_mux2_signals[0][10][29] , 
        \s_mux2_signals[0][10][28] , \s_mux2_signals[0][10][27] , 
        \s_mux2_signals[0][10][26] , \s_mux2_signals[0][10][25] , 
        \s_mux2_signals[0][10][24] , \s_mux2_signals[0][10][23] , 
        \s_mux2_signals[0][10][22] , \s_mux2_signals[0][10][21] , 
        \s_mux2_signals[0][10][20] , \s_mux2_signals[0][10][19] , 
        \s_mux2_signals[0][10][18] , \s_mux2_signals[0][10][17] , 
        \s_mux2_signals[0][10][16] , \s_mux2_signals[0][10][15] , 
        \s_mux2_signals[0][10][14] , \s_mux2_signals[0][10][13] , 
        \s_mux2_signals[0][10][12] , \s_mux2_signals[0][10][11] , 
        \s_mux2_signals[0][10][10] , \s_mux2_signals[0][10][9] , 
        \s_mux2_signals[0][10][8] , \s_mux2_signals[0][10][7] , 
        \s_mux2_signals[0][10][6] , \s_mux2_signals[0][10][5] , 
        \s_mux2_signals[0][10][4] , \s_mux2_signals[0][10][3] , 
        \s_mux2_signals[0][10][2] , \s_mux2_signals[0][10][1] , 
        \s_mux2_signals[0][10][0] }) );
  NRegister_N32_21 Ri_11 ( .clk(n9), .reset(n117), .data_in({n113, 
        RF_data_in[30:26], n105, n102, n99, RF_data_in[22], n95, n92, n89, n86, 
        n83, n80, n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, n44, 
        n41, n38, RF_data_in[1:0]}), .enable(n114), .load(
        s_load_Fdec_Tregs[11]), .data_out({\s_mux2_signals[0][11][31] , 
        \s_mux2_signals[0][11][30] , \s_mux2_signals[0][11][29] , 
        \s_mux2_signals[0][11][28] , \s_mux2_signals[0][11][27] , 
        \s_mux2_signals[0][11][26] , \s_mux2_signals[0][11][25] , 
        \s_mux2_signals[0][11][24] , \s_mux2_signals[0][11][23] , 
        \s_mux2_signals[0][11][22] , \s_mux2_signals[0][11][21] , 
        \s_mux2_signals[0][11][20] , \s_mux2_signals[0][11][19] , 
        \s_mux2_signals[0][11][18] , \s_mux2_signals[0][11][17] , 
        \s_mux2_signals[0][11][16] , \s_mux2_signals[0][11][15] , 
        \s_mux2_signals[0][11][14] , \s_mux2_signals[0][11][13] , 
        \s_mux2_signals[0][11][12] , \s_mux2_signals[0][11][11] , 
        \s_mux2_signals[0][11][10] , \s_mux2_signals[0][11][9] , 
        \s_mux2_signals[0][11][8] , \s_mux2_signals[0][11][7] , 
        \s_mux2_signals[0][11][6] , \s_mux2_signals[0][11][5] , 
        \s_mux2_signals[0][11][4] , \s_mux2_signals[0][11][3] , 
        \s_mux2_signals[0][11][2] , \s_mux2_signals[0][11][1] , 
        \s_mux2_signals[0][11][0] }) );
  NRegister_N32_20 Ri_12 ( .clk(n9), .reset(n117), .data_in({n113, 
        RF_data_in[30:26], n105, n102, n99, RF_data_in[22], n95, n92, n89, n86, 
        n83, n80, n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, n44, 
        n41, n38, RF_data_in[1:0]}), .enable(n114), .load(
        s_load_Fdec_Tregs[12]), .data_out({\s_mux2_signals[0][12][31] , 
        \s_mux2_signals[0][12][30] , \s_mux2_signals[0][12][29] , 
        \s_mux2_signals[0][12][28] , \s_mux2_signals[0][12][27] , 
        \s_mux2_signals[0][12][26] , \s_mux2_signals[0][12][25] , 
        \s_mux2_signals[0][12][24] , \s_mux2_signals[0][12][23] , 
        \s_mux2_signals[0][12][22] , \s_mux2_signals[0][12][21] , 
        \s_mux2_signals[0][12][20] , \s_mux2_signals[0][12][19] , 
        \s_mux2_signals[0][12][18] , \s_mux2_signals[0][12][17] , 
        \s_mux2_signals[0][12][16] , \s_mux2_signals[0][12][15] , 
        \s_mux2_signals[0][12][14] , \s_mux2_signals[0][12][13] , 
        \s_mux2_signals[0][12][12] , \s_mux2_signals[0][12][11] , 
        \s_mux2_signals[0][12][10] , \s_mux2_signals[0][12][9] , 
        \s_mux2_signals[0][12][8] , \s_mux2_signals[0][12][7] , 
        \s_mux2_signals[0][12][6] , \s_mux2_signals[0][12][5] , 
        \s_mux2_signals[0][12][4] , \s_mux2_signals[0][12][3] , 
        \s_mux2_signals[0][12][2] , \s_mux2_signals[0][12][1] , 
        \s_mux2_signals[0][12][0] }) );
  NRegister_N32_19 Ri_13 ( .clk(n9), .reset(n117), .data_in({n113, 
        RF_data_in[30:26], n105, n102, n99, RF_data_in[22], n95, n92, n89, n86, 
        n83, n80, n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, n44, 
        n41, n38, RF_data_in[1:0]}), .enable(n114), .load(
        s_load_Fdec_Tregs[13]), .data_out({\s_mux2_signals[0][13][31] , 
        \s_mux2_signals[0][13][30] , \s_mux2_signals[0][13][29] , 
        \s_mux2_signals[0][13][28] , \s_mux2_signals[0][13][27] , 
        \s_mux2_signals[0][13][26] , \s_mux2_signals[0][13][25] , 
        \s_mux2_signals[0][13][24] , \s_mux2_signals[0][13][23] , 
        \s_mux2_signals[0][13][22] , \s_mux2_signals[0][13][21] , 
        \s_mux2_signals[0][13][20] , \s_mux2_signals[0][13][19] , 
        \s_mux2_signals[0][13][18] , \s_mux2_signals[0][13][17] , 
        \s_mux2_signals[0][13][16] , \s_mux2_signals[0][13][15] , 
        \s_mux2_signals[0][13][14] , \s_mux2_signals[0][13][13] , 
        \s_mux2_signals[0][13][12] , \s_mux2_signals[0][13][11] , 
        \s_mux2_signals[0][13][10] , \s_mux2_signals[0][13][9] , 
        \s_mux2_signals[0][13][8] , \s_mux2_signals[0][13][7] , 
        \s_mux2_signals[0][13][6] , \s_mux2_signals[0][13][5] , 
        \s_mux2_signals[0][13][4] , \s_mux2_signals[0][13][3] , 
        \s_mux2_signals[0][13][2] , \s_mux2_signals[0][13][1] , 
        \s_mux2_signals[0][13][0] }) );
  NRegister_N32_18 Ri_14 ( .clk(n9), .reset(n117), .data_in({n113, 
        RF_data_in[30:26], n105, n102, n99, RF_data_in[22], n95, n92, n89, n86, 
        n83, n80, n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, n44, 
        n41, n38, RF_data_in[1:0]}), .enable(n114), .load(
        s_load_Fdec_Tregs[14]), .data_out({\s_mux2_signals[0][14][31] , 
        \s_mux2_signals[0][14][30] , \s_mux2_signals[0][14][29] , 
        \s_mux2_signals[0][14][28] , \s_mux2_signals[0][14][27] , 
        \s_mux2_signals[0][14][26] , \s_mux2_signals[0][14][25] , 
        \s_mux2_signals[0][14][24] , \s_mux2_signals[0][14][23] , 
        \s_mux2_signals[0][14][22] , \s_mux2_signals[0][14][21] , 
        \s_mux2_signals[0][14][20] , \s_mux2_signals[0][14][19] , 
        \s_mux2_signals[0][14][18] , \s_mux2_signals[0][14][17] , 
        \s_mux2_signals[0][14][16] , \s_mux2_signals[0][14][15] , 
        \s_mux2_signals[0][14][14] , \s_mux2_signals[0][14][13] , 
        \s_mux2_signals[0][14][12] , \s_mux2_signals[0][14][11] , 
        \s_mux2_signals[0][14][10] , \s_mux2_signals[0][14][9] , 
        \s_mux2_signals[0][14][8] , \s_mux2_signals[0][14][7] , 
        \s_mux2_signals[0][14][6] , \s_mux2_signals[0][14][5] , 
        \s_mux2_signals[0][14][4] , \s_mux2_signals[0][14][3] , 
        \s_mux2_signals[0][14][2] , \s_mux2_signals[0][14][1] , 
        \s_mux2_signals[0][14][0] }) );
  NRegister_N32_17 Ri_15 ( .clk(n9), .reset(n118), .data_in({RF_data_in[31:26], 
        n106, n103, n100, RF_data_in[22], n96, n93, n90, n87, n84, n81, n78, 
        n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, n39, 
        RF_data_in[1:0]}), .enable(n115), .load(s_load_Fdec_Tregs[15]), 
        .data_out({\s_mux2_signals[0][15][31] , \s_mux2_signals[0][15][30] , 
        \s_mux2_signals[0][15][29] , \s_mux2_signals[0][15][28] , 
        \s_mux2_signals[0][15][27] , \s_mux2_signals[0][15][26] , 
        \s_mux2_signals[0][15][25] , \s_mux2_signals[0][15][24] , 
        \s_mux2_signals[0][15][23] , \s_mux2_signals[0][15][22] , 
        \s_mux2_signals[0][15][21] , \s_mux2_signals[0][15][20] , 
        \s_mux2_signals[0][15][19] , \s_mux2_signals[0][15][18] , 
        \s_mux2_signals[0][15][17] , \s_mux2_signals[0][15][16] , 
        \s_mux2_signals[0][15][15] , \s_mux2_signals[0][15][14] , 
        \s_mux2_signals[0][15][13] , \s_mux2_signals[0][15][12] , 
        \s_mux2_signals[0][15][11] , \s_mux2_signals[0][15][10] , 
        \s_mux2_signals[0][15][9] , \s_mux2_signals[0][15][8] , 
        \s_mux2_signals[0][15][7] , \s_mux2_signals[0][15][6] , 
        \s_mux2_signals[0][15][5] , \s_mux2_signals[0][15][4] , 
        \s_mux2_signals[0][15][3] , \s_mux2_signals[0][15][2] , 
        \s_mux2_signals[0][15][1] , \s_mux2_signals[0][15][0] }) );
  NRegister_N32_16 Ri_16 ( .clk(n9), .reset(n118), .data_in({RF_data_in[31:26], 
        n106, n103, n100, RF_data_in[22], n96, n93, n90, n87, n84, n81, n78, 
        n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, n39, 
        RF_data_in[1:0]}), .enable(n115), .load(s_load_Fdec_Tregs[16]), 
        .data_out({\s_mux2_signals[0][16][31] , \s_mux2_signals[0][16][30] , 
        \s_mux2_signals[0][16][29] , \s_mux2_signals[0][16][28] , 
        \s_mux2_signals[0][16][27] , \s_mux2_signals[0][16][26] , 
        \s_mux2_signals[0][16][25] , \s_mux2_signals[0][16][24] , 
        \s_mux2_signals[0][16][23] , \s_mux2_signals[0][16][22] , 
        \s_mux2_signals[0][16][21] , \s_mux2_signals[0][16][20] , 
        \s_mux2_signals[0][16][19] , \s_mux2_signals[0][16][18] , 
        \s_mux2_signals[0][16][17] , \s_mux2_signals[0][16][16] , 
        \s_mux2_signals[0][16][15] , \s_mux2_signals[0][16][14] , 
        \s_mux2_signals[0][16][13] , \s_mux2_signals[0][16][12] , 
        \s_mux2_signals[0][16][11] , \s_mux2_signals[0][16][10] , 
        \s_mux2_signals[0][16][9] , \s_mux2_signals[0][16][8] , 
        \s_mux2_signals[0][16][7] , \s_mux2_signals[0][16][6] , 
        \s_mux2_signals[0][16][5] , \s_mux2_signals[0][16][4] , 
        \s_mux2_signals[0][16][3] , \s_mux2_signals[0][16][2] , 
        \s_mux2_signals[0][16][1] , \s_mux2_signals[0][16][0] }) );
  NRegister_N32_15 Ri_17 ( .clk(n9), .reset(n118), .data_in({RF_data_in[31:26], 
        n106, n103, n100, RF_data_in[22], n96, n93, n90, n87, n84, n81, n78, 
        n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, n39, 
        RF_data_in[1:0]}), .enable(n115), .load(s_load_Fdec_Tregs[17]), 
        .data_out({\s_mux2_signals[0][17][31] , \s_mux2_signals[0][17][30] , 
        \s_mux2_signals[0][17][29] , \s_mux2_signals[0][17][28] , 
        \s_mux2_signals[0][17][27] , \s_mux2_signals[0][17][26] , 
        \s_mux2_signals[0][17][25] , \s_mux2_signals[0][17][24] , 
        \s_mux2_signals[0][17][23] , \s_mux2_signals[0][17][22] , 
        \s_mux2_signals[0][17][21] , \s_mux2_signals[0][17][20] , 
        \s_mux2_signals[0][17][19] , \s_mux2_signals[0][17][18] , 
        \s_mux2_signals[0][17][17] , \s_mux2_signals[0][17][16] , 
        \s_mux2_signals[0][17][15] , \s_mux2_signals[0][17][14] , 
        \s_mux2_signals[0][17][13] , \s_mux2_signals[0][17][12] , 
        \s_mux2_signals[0][17][11] , \s_mux2_signals[0][17][10] , 
        \s_mux2_signals[0][17][9] , \s_mux2_signals[0][17][8] , 
        \s_mux2_signals[0][17][7] , \s_mux2_signals[0][17][6] , 
        \s_mux2_signals[0][17][5] , \s_mux2_signals[0][17][4] , 
        \s_mux2_signals[0][17][3] , \s_mux2_signals[0][17][2] , 
        \s_mux2_signals[0][17][1] , \s_mux2_signals[0][17][0] }) );
  NRegister_N32_14 Ri_18 ( .clk(n9), .reset(n119), .data_in({RF_data_in[31], 
        n112, n111, n110, n109, n108, n107, n104, n101, n98, n97, n94, n91, 
        n88, n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, 
        n46, n43, n40, n37, n36}), .enable(n116), .load(s_load_Fdec_Tregs[18]), 
        .data_out({\s_mux2_signals[0][18][31] , \s_mux2_signals[0][18][30] , 
        \s_mux2_signals[0][18][29] , \s_mux2_signals[0][18][28] , 
        \s_mux2_signals[0][18][27] , \s_mux2_signals[0][18][26] , 
        \s_mux2_signals[0][18][25] , \s_mux2_signals[0][18][24] , 
        \s_mux2_signals[0][18][23] , \s_mux2_signals[0][18][22] , 
        \s_mux2_signals[0][18][21] , \s_mux2_signals[0][18][20] , 
        \s_mux2_signals[0][18][19] , \s_mux2_signals[0][18][18] , 
        \s_mux2_signals[0][18][17] , \s_mux2_signals[0][18][16] , 
        \s_mux2_signals[0][18][15] , \s_mux2_signals[0][18][14] , 
        \s_mux2_signals[0][18][13] , \s_mux2_signals[0][18][12] , 
        \s_mux2_signals[0][18][11] , \s_mux2_signals[0][18][10] , 
        \s_mux2_signals[0][18][9] , \s_mux2_signals[0][18][8] , 
        \s_mux2_signals[0][18][7] , \s_mux2_signals[0][18][6] , 
        \s_mux2_signals[0][18][5] , \s_mux2_signals[0][18][4] , 
        \s_mux2_signals[0][18][3] , \s_mux2_signals[0][18][2] , 
        \s_mux2_signals[0][18][1] , \s_mux2_signals[0][18][0] }) );
  NRegister_N32_13 Ri_19 ( .clk(n9), .reset(n118), .data_in({RF_data_in[31:26], 
        n106, n103, n100, RF_data_in[22], n96, n93, n90, n87, n84, n81, n78, 
        n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, n39, 
        RF_data_in[1:0]}), .enable(n115), .load(s_load_Fdec_Tregs[19]), 
        .data_out({\s_mux2_signals[0][19][31] , \s_mux2_signals[0][19][30] , 
        \s_mux2_signals[0][19][29] , \s_mux2_signals[0][19][28] , 
        \s_mux2_signals[0][19][27] , \s_mux2_signals[0][19][26] , 
        \s_mux2_signals[0][19][25] , \s_mux2_signals[0][19][24] , 
        \s_mux2_signals[0][19][23] , \s_mux2_signals[0][19][22] , 
        \s_mux2_signals[0][19][21] , \s_mux2_signals[0][19][20] , 
        \s_mux2_signals[0][19][19] , \s_mux2_signals[0][19][18] , 
        \s_mux2_signals[0][19][17] , \s_mux2_signals[0][19][16] , 
        \s_mux2_signals[0][19][15] , \s_mux2_signals[0][19][14] , 
        \s_mux2_signals[0][19][13] , \s_mux2_signals[0][19][12] , 
        \s_mux2_signals[0][19][11] , \s_mux2_signals[0][19][10] , 
        \s_mux2_signals[0][19][9] , \s_mux2_signals[0][19][8] , 
        \s_mux2_signals[0][19][7] , \s_mux2_signals[0][19][6] , 
        \s_mux2_signals[0][19][5] , \s_mux2_signals[0][19][4] , 
        \s_mux2_signals[0][19][3] , \s_mux2_signals[0][19][2] , 
        \s_mux2_signals[0][19][1] , \s_mux2_signals[0][19][0] }) );
  NRegister_N32_12 Ri_20 ( .clk(n9), .reset(n118), .data_in({RF_data_in[31:26], 
        n106, n103, n100, RF_data_in[22], n96, n93, n90, n87, n84, n81, n78, 
        n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, n39, 
        RF_data_in[1:0]}), .enable(n115), .load(s_load_Fdec_Tregs[20]), 
        .data_out({\s_mux2_signals[0][20][31] , \s_mux2_signals[0][20][30] , 
        \s_mux2_signals[0][20][29] , \s_mux2_signals[0][20][28] , 
        \s_mux2_signals[0][20][27] , \s_mux2_signals[0][20][26] , 
        \s_mux2_signals[0][20][25] , \s_mux2_signals[0][20][24] , 
        \s_mux2_signals[0][20][23] , \s_mux2_signals[0][20][22] , 
        \s_mux2_signals[0][20][21] , \s_mux2_signals[0][20][20] , 
        \s_mux2_signals[0][20][19] , \s_mux2_signals[0][20][18] , 
        \s_mux2_signals[0][20][17] , \s_mux2_signals[0][20][16] , 
        \s_mux2_signals[0][20][15] , \s_mux2_signals[0][20][14] , 
        \s_mux2_signals[0][20][13] , \s_mux2_signals[0][20][12] , 
        \s_mux2_signals[0][20][11] , \s_mux2_signals[0][20][10] , 
        \s_mux2_signals[0][20][9] , \s_mux2_signals[0][20][8] , 
        \s_mux2_signals[0][20][7] , \s_mux2_signals[0][20][6] , 
        \s_mux2_signals[0][20][5] , \s_mux2_signals[0][20][4] , 
        \s_mux2_signals[0][20][3] , \s_mux2_signals[0][20][2] , 
        \s_mux2_signals[0][20][1] , \s_mux2_signals[0][20][0] }) );
  NRegister_N32_11 Ri_21 ( .clk(n9), .reset(n118), .data_in({RF_data_in[31:26], 
        n106, n103, n100, RF_data_in[22], n96, n93, n90, n87, n84, n81, n78, 
        n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, n39, 
        RF_data_in[1:0]}), .enable(n115), .load(s_load_Fdec_Tregs[21]), 
        .data_out({\s_mux2_signals[0][21][31] , \s_mux2_signals[0][21][30] , 
        \s_mux2_signals[0][21][29] , \s_mux2_signals[0][21][28] , 
        \s_mux2_signals[0][21][27] , \s_mux2_signals[0][21][26] , 
        \s_mux2_signals[0][21][25] , \s_mux2_signals[0][21][24] , 
        \s_mux2_signals[0][21][23] , \s_mux2_signals[0][21][22] , 
        \s_mux2_signals[0][21][21] , \s_mux2_signals[0][21][20] , 
        \s_mux2_signals[0][21][19] , \s_mux2_signals[0][21][18] , 
        \s_mux2_signals[0][21][17] , \s_mux2_signals[0][21][16] , 
        \s_mux2_signals[0][21][15] , \s_mux2_signals[0][21][14] , 
        \s_mux2_signals[0][21][13] , \s_mux2_signals[0][21][12] , 
        \s_mux2_signals[0][21][11] , \s_mux2_signals[0][21][10] , 
        \s_mux2_signals[0][21][9] , \s_mux2_signals[0][21][8] , 
        \s_mux2_signals[0][21][7] , \s_mux2_signals[0][21][6] , 
        \s_mux2_signals[0][21][5] , \s_mux2_signals[0][21][4] , 
        \s_mux2_signals[0][21][3] , \s_mux2_signals[0][21][2] , 
        \s_mux2_signals[0][21][1] , \s_mux2_signals[0][21][0] }) );
  NRegister_N32_10 Ri_22 ( .clk(n9), .reset(n118), .data_in({RF_data_in[31:26], 
        n106, n103, n100, RF_data_in[22], n96, n93, n90, n87, n84, n81, n78, 
        n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, n39, 
        RF_data_in[1:0]}), .enable(n115), .load(s_load_Fdec_Tregs[22]), 
        .data_out({\s_mux2_signals[0][22][31] , \s_mux2_signals[0][22][30] , 
        \s_mux2_signals[0][22][29] , \s_mux2_signals[0][22][28] , 
        \s_mux2_signals[0][22][27] , \s_mux2_signals[0][22][26] , 
        \s_mux2_signals[0][22][25] , \s_mux2_signals[0][22][24] , 
        \s_mux2_signals[0][22][23] , \s_mux2_signals[0][22][22] , 
        \s_mux2_signals[0][22][21] , \s_mux2_signals[0][22][20] , 
        \s_mux2_signals[0][22][19] , \s_mux2_signals[0][22][18] , 
        \s_mux2_signals[0][22][17] , \s_mux2_signals[0][22][16] , 
        \s_mux2_signals[0][22][15] , \s_mux2_signals[0][22][14] , 
        \s_mux2_signals[0][22][13] , \s_mux2_signals[0][22][12] , 
        \s_mux2_signals[0][22][11] , \s_mux2_signals[0][22][10] , 
        \s_mux2_signals[0][22][9] , \s_mux2_signals[0][22][8] , 
        \s_mux2_signals[0][22][7] , \s_mux2_signals[0][22][6] , 
        \s_mux2_signals[0][22][5] , \s_mux2_signals[0][22][4] , 
        \s_mux2_signals[0][22][3] , \s_mux2_signals[0][22][2] , 
        \s_mux2_signals[0][22][1] , \s_mux2_signals[0][22][0] }) );
  NRegister_N32_9 Ri_23 ( .clk(n9), .reset(n118), .data_in({RF_data_in[31:26], 
        n106, n103, n100, RF_data_in[22], n96, n93, n90, n87, n84, n81, n78, 
        n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, n39, 
        RF_data_in[1:0]}), .enable(n115), .load(s_load_Fdec_Tregs[23]), 
        .data_out({\s_mux2_signals[0][23][31] , \s_mux2_signals[0][23][30] , 
        \s_mux2_signals[0][23][29] , \s_mux2_signals[0][23][28] , 
        \s_mux2_signals[0][23][27] , \s_mux2_signals[0][23][26] , 
        \s_mux2_signals[0][23][25] , \s_mux2_signals[0][23][24] , 
        \s_mux2_signals[0][23][23] , \s_mux2_signals[0][23][22] , 
        \s_mux2_signals[0][23][21] , \s_mux2_signals[0][23][20] , 
        \s_mux2_signals[0][23][19] , \s_mux2_signals[0][23][18] , 
        \s_mux2_signals[0][23][17] , \s_mux2_signals[0][23][16] , 
        \s_mux2_signals[0][23][15] , \s_mux2_signals[0][23][14] , 
        \s_mux2_signals[0][23][13] , \s_mux2_signals[0][23][12] , 
        \s_mux2_signals[0][23][11] , \s_mux2_signals[0][23][10] , 
        \s_mux2_signals[0][23][9] , \s_mux2_signals[0][23][8] , 
        \s_mux2_signals[0][23][7] , \s_mux2_signals[0][23][6] , 
        \s_mux2_signals[0][23][5] , \s_mux2_signals[0][23][4] , 
        \s_mux2_signals[0][23][3] , \s_mux2_signals[0][23][2] , 
        \s_mux2_signals[0][23][1] , \s_mux2_signals[0][23][0] }) );
  NRegister_N32_8 Ri_24 ( .clk(n9), .reset(n118), .data_in({RF_data_in[31:26], 
        n106, n103, n100, RF_data_in[22], n96, n93, n90, n87, n84, n81, n78, 
        n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, n39, 
        RF_data_in[1:0]}), .enable(n115), .load(s_load_Fdec_Tregs[24]), 
        .data_out({\s_mux2_signals[0][24][31] , \s_mux2_signals[0][24][30] , 
        \s_mux2_signals[0][24][29] , \s_mux2_signals[0][24][28] , 
        \s_mux2_signals[0][24][27] , \s_mux2_signals[0][24][26] , 
        \s_mux2_signals[0][24][25] , \s_mux2_signals[0][24][24] , 
        \s_mux2_signals[0][24][23] , \s_mux2_signals[0][24][22] , 
        \s_mux2_signals[0][24][21] , \s_mux2_signals[0][24][20] , 
        \s_mux2_signals[0][24][19] , \s_mux2_signals[0][24][18] , 
        \s_mux2_signals[0][24][17] , \s_mux2_signals[0][24][16] , 
        \s_mux2_signals[0][24][15] , \s_mux2_signals[0][24][14] , 
        \s_mux2_signals[0][24][13] , \s_mux2_signals[0][24][12] , 
        \s_mux2_signals[0][24][11] , \s_mux2_signals[0][24][10] , 
        \s_mux2_signals[0][24][9] , \s_mux2_signals[0][24][8] , 
        \s_mux2_signals[0][24][7] , \s_mux2_signals[0][24][6] , 
        \s_mux2_signals[0][24][5] , \s_mux2_signals[0][24][4] , 
        \s_mux2_signals[0][24][3] , \s_mux2_signals[0][24][2] , 
        \s_mux2_signals[0][24][1] , \s_mux2_signals[0][24][0] }) );
  NRegister_N32_7 Ri_25 ( .clk(n9), .reset(n118), .data_in({RF_data_in[31:26], 
        n106, n103, n100, RF_data_in[22], n96, n93, n90, n87, n84, n81, n78, 
        n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, n39, 
        RF_data_in[1:0]}), .enable(n115), .load(s_load_Fdec_Tregs[25]), 
        .data_out({\s_mux2_signals[0][25][31] , \s_mux2_signals[0][25][30] , 
        \s_mux2_signals[0][25][29] , \s_mux2_signals[0][25][28] , 
        \s_mux2_signals[0][25][27] , \s_mux2_signals[0][25][26] , 
        \s_mux2_signals[0][25][25] , \s_mux2_signals[0][25][24] , 
        \s_mux2_signals[0][25][23] , \s_mux2_signals[0][25][22] , 
        \s_mux2_signals[0][25][21] , \s_mux2_signals[0][25][20] , 
        \s_mux2_signals[0][25][19] , \s_mux2_signals[0][25][18] , 
        \s_mux2_signals[0][25][17] , \s_mux2_signals[0][25][16] , 
        \s_mux2_signals[0][25][15] , \s_mux2_signals[0][25][14] , 
        \s_mux2_signals[0][25][13] , \s_mux2_signals[0][25][12] , 
        \s_mux2_signals[0][25][11] , \s_mux2_signals[0][25][10] , 
        \s_mux2_signals[0][25][9] , \s_mux2_signals[0][25][8] , 
        \s_mux2_signals[0][25][7] , \s_mux2_signals[0][25][6] , 
        \s_mux2_signals[0][25][5] , \s_mux2_signals[0][25][4] , 
        \s_mux2_signals[0][25][3] , \s_mux2_signals[0][25][2] , 
        \s_mux2_signals[0][25][1] , \s_mux2_signals[0][25][0] }) );
  NRegister_N32_6 Ri_26 ( .clk(n9), .reset(n118), .data_in({RF_data_in[31:26], 
        n106, n103, n100, RF_data_in[22], n96, n93, n90, n87, n84, n81, n78, 
        n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, n39, 
        RF_data_in[1:0]}), .enable(n115), .load(s_load_Fdec_Tregs[26]), 
        .data_out({\s_mux2_signals[0][26][31] , \s_mux2_signals[0][26][30] , 
        \s_mux2_signals[0][26][29] , \s_mux2_signals[0][26][28] , 
        \s_mux2_signals[0][26][27] , \s_mux2_signals[0][26][26] , 
        \s_mux2_signals[0][26][25] , \s_mux2_signals[0][26][24] , 
        \s_mux2_signals[0][26][23] , \s_mux2_signals[0][26][22] , 
        \s_mux2_signals[0][26][21] , \s_mux2_signals[0][26][20] , 
        \s_mux2_signals[0][26][19] , \s_mux2_signals[0][26][18] , 
        \s_mux2_signals[0][26][17] , \s_mux2_signals[0][26][16] , 
        \s_mux2_signals[0][26][15] , \s_mux2_signals[0][26][14] , 
        \s_mux2_signals[0][26][13] , \s_mux2_signals[0][26][12] , 
        \s_mux2_signals[0][26][11] , \s_mux2_signals[0][26][10] , 
        \s_mux2_signals[0][26][9] , \s_mux2_signals[0][26][8] , 
        \s_mux2_signals[0][26][7] , \s_mux2_signals[0][26][6] , 
        \s_mux2_signals[0][26][5] , \s_mux2_signals[0][26][4] , 
        \s_mux2_signals[0][26][3] , \s_mux2_signals[0][26][2] , 
        \s_mux2_signals[0][26][1] , \s_mux2_signals[0][26][0] }) );
  NRegister_N32_5 Ri_27 ( .clk(n9), .reset(n119), .data_in({RF_data_in[31], 
        n112, n111, n110, n109, n108, n107, n104, n101, n98, n97, n94, n91, 
        n88, n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, 
        n46, n43, n40, n37, n36}), .enable(n116), .load(s_load_Fdec_Tregs[27]), 
        .data_out({\s_mux2_signals[0][27][31] , \s_mux2_signals[0][27][30] , 
        \s_mux2_signals[0][27][29] , \s_mux2_signals[0][27][28] , 
        \s_mux2_signals[0][27][27] , \s_mux2_signals[0][27][26] , 
        \s_mux2_signals[0][27][25] , \s_mux2_signals[0][27][24] , 
        \s_mux2_signals[0][27][23] , \s_mux2_signals[0][27][22] , 
        \s_mux2_signals[0][27][21] , \s_mux2_signals[0][27][20] , 
        \s_mux2_signals[0][27][19] , \s_mux2_signals[0][27][18] , 
        \s_mux2_signals[0][27][17] , \s_mux2_signals[0][27][16] , 
        \s_mux2_signals[0][27][15] , \s_mux2_signals[0][27][14] , 
        \s_mux2_signals[0][27][13] , \s_mux2_signals[0][27][12] , 
        \s_mux2_signals[0][27][11] , \s_mux2_signals[0][27][10] , 
        \s_mux2_signals[0][27][9] , \s_mux2_signals[0][27][8] , 
        \s_mux2_signals[0][27][7] , \s_mux2_signals[0][27][6] , 
        \s_mux2_signals[0][27][5] , \s_mux2_signals[0][27][4] , 
        \s_mux2_signals[0][27][3] , \s_mux2_signals[0][27][2] , 
        \s_mux2_signals[0][27][1] , \s_mux2_signals[0][27][0] }) );
  NRegister_N32_4 Ri_28 ( .clk(n9), .reset(n118), .data_in({RF_data_in[31:26], 
        n106, n103, n100, RF_data_in[22], n96, n93, n90, n87, n84, n81, n78, 
        n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, n39, 
        RF_data_in[1:0]}), .enable(n115), .load(s_load_Fdec_Tregs[28]), 
        .data_out({\s_mux2_signals[0][28][31] , \s_mux2_signals[0][28][30] , 
        \s_mux2_signals[0][28][29] , \s_mux2_signals[0][28][28] , 
        \s_mux2_signals[0][28][27] , \s_mux2_signals[0][28][26] , 
        \s_mux2_signals[0][28][25] , \s_mux2_signals[0][28][24] , 
        \s_mux2_signals[0][28][23] , \s_mux2_signals[0][28][22] , 
        \s_mux2_signals[0][28][21] , \s_mux2_signals[0][28][20] , 
        \s_mux2_signals[0][28][19] , \s_mux2_signals[0][28][18] , 
        \s_mux2_signals[0][28][17] , \s_mux2_signals[0][28][16] , 
        \s_mux2_signals[0][28][15] , \s_mux2_signals[0][28][14] , 
        \s_mux2_signals[0][28][13] , \s_mux2_signals[0][28][12] , 
        \s_mux2_signals[0][28][11] , \s_mux2_signals[0][28][10] , 
        \s_mux2_signals[0][28][9] , \s_mux2_signals[0][28][8] , 
        \s_mux2_signals[0][28][7] , \s_mux2_signals[0][28][6] , 
        \s_mux2_signals[0][28][5] , \s_mux2_signals[0][28][4] , 
        \s_mux2_signals[0][28][3] , \s_mux2_signals[0][28][2] , 
        \s_mux2_signals[0][28][1] , \s_mux2_signals[0][28][0] }) );
  NRegister_N32_3 Ri_29 ( .clk(n9), .reset(n119), .data_in({RF_data_in[31], 
        n112, n111, n110, n109, n108, n107, n104, n101, n98, n97, n94, n91, 
        n88, n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, 
        n46, n43, n40, n37, n36}), .enable(n116), .load(s_load_Fdec_Tregs[29]), 
        .data_out({\s_mux2_signals[0][29][31] , \s_mux2_signals[0][29][30] , 
        \s_mux2_signals[0][29][29] , \s_mux2_signals[0][29][28] , 
        \s_mux2_signals[0][29][27] , \s_mux2_signals[0][29][26] , 
        \s_mux2_signals[0][29][25] , \s_mux2_signals[0][29][24] , 
        \s_mux2_signals[0][29][23] , \s_mux2_signals[0][29][22] , 
        \s_mux2_signals[0][29][21] , \s_mux2_signals[0][29][20] , 
        \s_mux2_signals[0][29][19] , \s_mux2_signals[0][29][18] , 
        \s_mux2_signals[0][29][17] , \s_mux2_signals[0][29][16] , 
        \s_mux2_signals[0][29][15] , \s_mux2_signals[0][29][14] , 
        \s_mux2_signals[0][29][13] , \s_mux2_signals[0][29][12] , 
        \s_mux2_signals[0][29][11] , \s_mux2_signals[0][29][10] , 
        \s_mux2_signals[0][29][9] , \s_mux2_signals[0][29][8] , 
        \s_mux2_signals[0][29][7] , \s_mux2_signals[0][29][6] , 
        \s_mux2_signals[0][29][5] , \s_mux2_signals[0][29][4] , 
        \s_mux2_signals[0][29][3] , \s_mux2_signals[0][29][2] , 
        \s_mux2_signals[0][29][1] , \s_mux2_signals[0][29][0] }) );
  NRegister_N32_2 Ri_30 ( .clk(n9), .reset(n119), .data_in({RF_data_in[31], 
        n112, n111, n110, n109, n108, n107, n104, n101, n98, n97, n94, n91, 
        n88, n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, 
        n46, n43, n40, n37, n36}), .enable(n116), .load(s_load_Fdec_Tregs[30]), 
        .data_out({\s_mux2_signals[0][30][31] , \s_mux2_signals[0][30][30] , 
        \s_mux2_signals[0][30][29] , \s_mux2_signals[0][30][28] , 
        \s_mux2_signals[0][30][27] , \s_mux2_signals[0][30][26] , 
        \s_mux2_signals[0][30][25] , \s_mux2_signals[0][30][24] , 
        \s_mux2_signals[0][30][23] , \s_mux2_signals[0][30][22] , 
        \s_mux2_signals[0][30][21] , \s_mux2_signals[0][30][20] , 
        \s_mux2_signals[0][30][19] , \s_mux2_signals[0][30][18] , 
        \s_mux2_signals[0][30][17] , \s_mux2_signals[0][30][16] , 
        \s_mux2_signals[0][30][15] , \s_mux2_signals[0][30][14] , 
        \s_mux2_signals[0][30][13] , \s_mux2_signals[0][30][12] , 
        \s_mux2_signals[0][30][11] , \s_mux2_signals[0][30][10] , 
        \s_mux2_signals[0][30][9] , \s_mux2_signals[0][30][8] , 
        \s_mux2_signals[0][30][7] , \s_mux2_signals[0][30][6] , 
        \s_mux2_signals[0][30][5] , \s_mux2_signals[0][30][4] , 
        \s_mux2_signals[0][30][3] , \s_mux2_signals[0][30][2] , 
        \s_mux2_signals[0][30][1] , \s_mux2_signals[0][30][0] }) );
  NRegister_N32_1 Ri_31 ( .clk(n9), .reset(n119), .data_in({RF_data_in[31], 
        n112, n111, n110, n109, n108, n107, n104, n101, n98, n97, n94, n91, 
        n88, n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, 
        n46, n43, n40, n37, n36}), .enable(n116), .load(s_load_Fdec_Tregs[31]), 
        .data_out({\s_mux2_signals[0][31][31] , \s_mux2_signals[0][31][30] , 
        \s_mux2_signals[0][31][29] , \s_mux2_signals[0][31][28] , 
        \s_mux2_signals[0][31][27] , \s_mux2_signals[0][31][26] , 
        \s_mux2_signals[0][31][25] , \s_mux2_signals[0][31][24] , 
        \s_mux2_signals[0][31][23] , \s_mux2_signals[0][31][22] , 
        \s_mux2_signals[0][31][21] , \s_mux2_signals[0][31][20] , 
        \s_mux2_signals[0][31][19] , \s_mux2_signals[0][31][18] , 
        \s_mux2_signals[0][31][17] , \s_mux2_signals[0][31][16] , 
        \s_mux2_signals[0][31][15] , \s_mux2_signals[0][31][14] , 
        \s_mux2_signals[0][31][13] , \s_mux2_signals[0][31][12] , 
        \s_mux2_signals[0][31][11] , \s_mux2_signals[0][31][10] , 
        \s_mux2_signals[0][31][9] , \s_mux2_signals[0][31][8] , 
        \s_mux2_signals[0][31][7] , \s_mux2_signals[0][31][6] , 
        \s_mux2_signals[0][31][5] , \s_mux2_signals[0][31][4] , 
        \s_mux2_signals[0][31][3] , \s_mux2_signals[0][31][2] , 
        \s_mux2_signals[0][31][1] , \s_mux2_signals[0][31][0] }) );
  Mux_NBit_2x1_NBIT_IN32_79 MUX1_0_0 ( .port0({\s_mux2_signals[0][0][31] , 
        \s_mux2_signals[0][0][30] , \s_mux2_signals[0][0][29] , 
        \s_mux2_signals[0][0][28] , \s_mux2_signals[0][0][27] , 
        \s_mux2_signals[0][0][26] , \s_mux2_signals[0][0][25] , 
        \s_mux2_signals[0][0][24] , \s_mux2_signals[0][0][23] , 
        \s_mux2_signals[0][0][22] , \s_mux2_signals[0][0][21] , 
        \s_mux2_signals[0][0][20] , \s_mux2_signals[0][0][19] , 
        \s_mux2_signals[0][0][18] , \s_mux2_signals[0][0][17] , 
        \s_mux2_signals[0][0][16] , \s_mux2_signals[0][0][15] , 
        \s_mux2_signals[0][0][14] , \s_mux2_signals[0][0][13] , 
        \s_mux2_signals[0][0][12] , \s_mux2_signals[0][0][11] , 
        \s_mux2_signals[0][0][10] , \s_mux2_signals[0][0][9] , 
        \s_mux2_signals[0][0][8] , \s_mux2_signals[0][0][7] , 
        \s_mux2_signals[0][0][6] , \s_mux2_signals[0][0][5] , 
        \s_mux2_signals[0][0][4] , \s_mux2_signals[0][0][3] , 
        \s_mux2_signals[0][0][2] , \s_mux2_signals[0][0][1] , 
        \s_mux2_signals[0][0][0] }), .port1({\s_mux2_signals[0][1][31] , 
        \s_mux2_signals[0][1][30] , \s_mux2_signals[0][1][29] , 
        \s_mux2_signals[0][1][28] , \s_mux2_signals[0][1][27] , 
        \s_mux2_signals[0][1][26] , \s_mux2_signals[0][1][25] , 
        \s_mux2_signals[0][1][24] , \s_mux2_signals[0][1][23] , 
        \s_mux2_signals[0][1][22] , \s_mux2_signals[0][1][21] , 
        \s_mux2_signals[0][1][20] , \s_mux2_signals[0][1][19] , 
        \s_mux2_signals[0][1][18] , \s_mux2_signals[0][1][17] , 
        \s_mux2_signals[0][1][16] , \s_mux2_signals[0][1][15] , 
        \s_mux2_signals[0][1][14] , \s_mux2_signals[0][1][13] , 
        \s_mux2_signals[0][1][12] , \s_mux2_signals[0][1][11] , 
        \s_mux2_signals[0][1][10] , \s_mux2_signals[0][1][9] , 
        \s_mux2_signals[0][1][8] , \s_mux2_signals[0][1][7] , 
        \s_mux2_signals[0][1][6] , \s_mux2_signals[0][1][5] , 
        \s_mux2_signals[0][1][4] , \s_mux2_signals[0][1][3] , 
        \s_mux2_signals[0][1][2] , \s_mux2_signals[0][1][1] , 
        \s_mux2_signals[0][1][0] }), .sel(n24), .portY({
        \s_mux1_signals[1][0][31] , \s_mux1_signals[1][0][30] , 
        \s_mux1_signals[1][0][29] , \s_mux1_signals[1][0][28] , 
        \s_mux1_signals[1][0][27] , \s_mux1_signals[1][0][26] , 
        \s_mux1_signals[1][0][25] , \s_mux1_signals[1][0][24] , 
        \s_mux1_signals[1][0][23] , \s_mux1_signals[1][0][22] , 
        \s_mux1_signals[1][0][21] , \s_mux1_signals[1][0][20] , 
        \s_mux1_signals[1][0][19] , \s_mux1_signals[1][0][18] , 
        \s_mux1_signals[1][0][17] , \s_mux1_signals[1][0][16] , 
        \s_mux1_signals[1][0][15] , \s_mux1_signals[1][0][14] , 
        \s_mux1_signals[1][0][13] , \s_mux1_signals[1][0][12] , 
        \s_mux1_signals[1][0][11] , \s_mux1_signals[1][0][10] , 
        \s_mux1_signals[1][0][9] , \s_mux1_signals[1][0][8] , 
        \s_mux1_signals[1][0][7] , \s_mux1_signals[1][0][6] , 
        \s_mux1_signals[1][0][5] , \s_mux1_signals[1][0][4] , 
        \s_mux1_signals[1][0][3] , \s_mux1_signals[1][0][2] , 
        \s_mux1_signals[1][0][1] , \s_mux1_signals[1][0][0] }) );
  Mux_NBit_2x1_NBIT_IN32_78 MUX1_0_2 ( .port0({\s_mux2_signals[0][2][31] , 
        \s_mux2_signals[0][2][30] , \s_mux2_signals[0][2][29] , 
        \s_mux2_signals[0][2][28] , \s_mux2_signals[0][2][27] , 
        \s_mux2_signals[0][2][26] , \s_mux2_signals[0][2][25] , 
        \s_mux2_signals[0][2][24] , \s_mux2_signals[0][2][23] , 
        \s_mux2_signals[0][2][22] , \s_mux2_signals[0][2][21] , 
        \s_mux2_signals[0][2][20] , \s_mux2_signals[0][2][19] , 
        \s_mux2_signals[0][2][18] , \s_mux2_signals[0][2][17] , 
        \s_mux2_signals[0][2][16] , \s_mux2_signals[0][2][15] , 
        \s_mux2_signals[0][2][14] , \s_mux2_signals[0][2][13] , 
        \s_mux2_signals[0][2][12] , \s_mux2_signals[0][2][11] , 
        \s_mux2_signals[0][2][10] , \s_mux2_signals[0][2][9] , 
        \s_mux2_signals[0][2][8] , \s_mux2_signals[0][2][7] , 
        \s_mux2_signals[0][2][6] , \s_mux2_signals[0][2][5] , 
        \s_mux2_signals[0][2][4] , \s_mux2_signals[0][2][3] , 
        \s_mux2_signals[0][2][2] , \s_mux2_signals[0][2][1] , 
        \s_mux2_signals[0][2][0] }), .port1({\s_mux2_signals[0][3][31] , 
        \s_mux2_signals[0][3][30] , \s_mux2_signals[0][3][29] , 
        \s_mux2_signals[0][3][28] , \s_mux2_signals[0][3][27] , 
        \s_mux2_signals[0][3][26] , \s_mux2_signals[0][3][25] , 
        \s_mux2_signals[0][3][24] , \s_mux2_signals[0][3][23] , 
        \s_mux2_signals[0][3][22] , \s_mux2_signals[0][3][21] , 
        \s_mux2_signals[0][3][20] , \s_mux2_signals[0][3][19] , 
        \s_mux2_signals[0][3][18] , \s_mux2_signals[0][3][17] , 
        \s_mux2_signals[0][3][16] , \s_mux2_signals[0][3][15] , 
        \s_mux2_signals[0][3][14] , \s_mux2_signals[0][3][13] , 
        \s_mux2_signals[0][3][12] , \s_mux2_signals[0][3][11] , 
        \s_mux2_signals[0][3][10] , \s_mux2_signals[0][3][9] , 
        \s_mux2_signals[0][3][8] , \s_mux2_signals[0][3][7] , 
        \s_mux2_signals[0][3][6] , \s_mux2_signals[0][3][5] , 
        \s_mux2_signals[0][3][4] , \s_mux2_signals[0][3][3] , 
        \s_mux2_signals[0][3][2] , \s_mux2_signals[0][3][1] , 
        \s_mux2_signals[0][3][0] }), .sel(n22), .portY({
        \s_mux1_signals[1][2][31] , \s_mux1_signals[1][2][30] , 
        \s_mux1_signals[1][2][29] , \s_mux1_signals[1][2][28] , 
        \s_mux1_signals[1][2][27] , \s_mux1_signals[1][2][26] , 
        \s_mux1_signals[1][2][25] , \s_mux1_signals[1][2][24] , 
        \s_mux1_signals[1][2][23] , \s_mux1_signals[1][2][22] , 
        \s_mux1_signals[1][2][21] , \s_mux1_signals[1][2][20] , 
        \s_mux1_signals[1][2][19] , \s_mux1_signals[1][2][18] , 
        \s_mux1_signals[1][2][17] , \s_mux1_signals[1][2][16] , 
        \s_mux1_signals[1][2][15] , \s_mux1_signals[1][2][14] , 
        \s_mux1_signals[1][2][13] , \s_mux1_signals[1][2][12] , 
        \s_mux1_signals[1][2][11] , \s_mux1_signals[1][2][10] , 
        \s_mux1_signals[1][2][9] , \s_mux1_signals[1][2][8] , 
        \s_mux1_signals[1][2][7] , \s_mux1_signals[1][2][6] , 
        \s_mux1_signals[1][2][5] , \s_mux1_signals[1][2][4] , 
        \s_mux1_signals[1][2][3] , \s_mux1_signals[1][2][2] , 
        \s_mux1_signals[1][2][1] , \s_mux1_signals[1][2][0] }) );
  Mux_NBit_2x1_NBIT_IN32_77 MUX1_0_4 ( .port0({\s_mux2_signals[0][4][31] , 
        \s_mux2_signals[0][4][30] , \s_mux2_signals[0][4][29] , 
        \s_mux2_signals[0][4][28] , \s_mux2_signals[0][4][27] , 
        \s_mux2_signals[0][4][26] , \s_mux2_signals[0][4][25] , 
        \s_mux2_signals[0][4][24] , \s_mux2_signals[0][4][23] , 
        \s_mux2_signals[0][4][22] , \s_mux2_signals[0][4][21] , 
        \s_mux2_signals[0][4][20] , \s_mux2_signals[0][4][19] , 
        \s_mux2_signals[0][4][18] , \s_mux2_signals[0][4][17] , 
        \s_mux2_signals[0][4][16] , \s_mux2_signals[0][4][15] , 
        \s_mux2_signals[0][4][14] , \s_mux2_signals[0][4][13] , 
        \s_mux2_signals[0][4][12] , \s_mux2_signals[0][4][11] , 
        \s_mux2_signals[0][4][10] , \s_mux2_signals[0][4][9] , 
        \s_mux2_signals[0][4][8] , \s_mux2_signals[0][4][7] , 
        \s_mux2_signals[0][4][6] , \s_mux2_signals[0][4][5] , 
        \s_mux2_signals[0][4][4] , \s_mux2_signals[0][4][3] , 
        \s_mux2_signals[0][4][2] , \s_mux2_signals[0][4][1] , 
        \s_mux2_signals[0][4][0] }), .port1({\s_mux2_signals[0][5][31] , 
        \s_mux2_signals[0][5][30] , \s_mux2_signals[0][5][29] , 
        \s_mux2_signals[0][5][28] , \s_mux2_signals[0][5][27] , 
        \s_mux2_signals[0][5][26] , \s_mux2_signals[0][5][25] , 
        \s_mux2_signals[0][5][24] , \s_mux2_signals[0][5][23] , 
        \s_mux2_signals[0][5][22] , \s_mux2_signals[0][5][21] , 
        \s_mux2_signals[0][5][20] , \s_mux2_signals[0][5][19] , 
        \s_mux2_signals[0][5][18] , \s_mux2_signals[0][5][17] , 
        \s_mux2_signals[0][5][16] , \s_mux2_signals[0][5][15] , 
        \s_mux2_signals[0][5][14] , \s_mux2_signals[0][5][13] , 
        \s_mux2_signals[0][5][12] , \s_mux2_signals[0][5][11] , 
        \s_mux2_signals[0][5][10] , \s_mux2_signals[0][5][9] , 
        \s_mux2_signals[0][5][8] , \s_mux2_signals[0][5][7] , 
        \s_mux2_signals[0][5][6] , \s_mux2_signals[0][5][5] , 
        \s_mux2_signals[0][5][4] , \s_mux2_signals[0][5][3] , 
        \s_mux2_signals[0][5][2] , \s_mux2_signals[0][5][1] , 
        \s_mux2_signals[0][5][0] }), .sel(n22), .portY({
        \s_mux1_signals[1][4][31] , \s_mux1_signals[1][4][30] , 
        \s_mux1_signals[1][4][29] , \s_mux1_signals[1][4][28] , 
        \s_mux1_signals[1][4][27] , \s_mux1_signals[1][4][26] , 
        \s_mux1_signals[1][4][25] , \s_mux1_signals[1][4][24] , 
        \s_mux1_signals[1][4][23] , \s_mux1_signals[1][4][22] , 
        \s_mux1_signals[1][4][21] , \s_mux1_signals[1][4][20] , 
        \s_mux1_signals[1][4][19] , \s_mux1_signals[1][4][18] , 
        \s_mux1_signals[1][4][17] , \s_mux1_signals[1][4][16] , 
        \s_mux1_signals[1][4][15] , \s_mux1_signals[1][4][14] , 
        \s_mux1_signals[1][4][13] , \s_mux1_signals[1][4][12] , 
        \s_mux1_signals[1][4][11] , \s_mux1_signals[1][4][10] , 
        \s_mux1_signals[1][4][9] , \s_mux1_signals[1][4][8] , 
        \s_mux1_signals[1][4][7] , \s_mux1_signals[1][4][6] , 
        \s_mux1_signals[1][4][5] , \s_mux1_signals[1][4][4] , 
        \s_mux1_signals[1][4][3] , \s_mux1_signals[1][4][2] , 
        \s_mux1_signals[1][4][1] , \s_mux1_signals[1][4][0] }) );
  Mux_NBit_2x1_NBIT_IN32_76 MUX1_0_6 ( .port0({\s_mux2_signals[0][6][31] , 
        \s_mux2_signals[0][6][30] , \s_mux2_signals[0][6][29] , 
        \s_mux2_signals[0][6][28] , \s_mux2_signals[0][6][27] , 
        \s_mux2_signals[0][6][26] , \s_mux2_signals[0][6][25] , 
        \s_mux2_signals[0][6][24] , \s_mux2_signals[0][6][23] , 
        \s_mux2_signals[0][6][22] , \s_mux2_signals[0][6][21] , 
        \s_mux2_signals[0][6][20] , \s_mux2_signals[0][6][19] , 
        \s_mux2_signals[0][6][18] , \s_mux2_signals[0][6][17] , 
        \s_mux2_signals[0][6][16] , \s_mux2_signals[0][6][15] , 
        \s_mux2_signals[0][6][14] , \s_mux2_signals[0][6][13] , 
        \s_mux2_signals[0][6][12] , \s_mux2_signals[0][6][11] , 
        \s_mux2_signals[0][6][10] , \s_mux2_signals[0][6][9] , 
        \s_mux2_signals[0][6][8] , \s_mux2_signals[0][6][7] , 
        \s_mux2_signals[0][6][6] , \s_mux2_signals[0][6][5] , 
        \s_mux2_signals[0][6][4] , \s_mux2_signals[0][6][3] , 
        \s_mux2_signals[0][6][2] , \s_mux2_signals[0][6][1] , 
        \s_mux2_signals[0][6][0] }), .port1({\s_mux2_signals[0][7][31] , 
        \s_mux2_signals[0][7][30] , \s_mux2_signals[0][7][29] , 
        \s_mux2_signals[0][7][28] , \s_mux2_signals[0][7][27] , 
        \s_mux2_signals[0][7][26] , \s_mux2_signals[0][7][25] , 
        \s_mux2_signals[0][7][24] , \s_mux2_signals[0][7][23] , 
        \s_mux2_signals[0][7][22] , \s_mux2_signals[0][7][21] , 
        \s_mux2_signals[0][7][20] , \s_mux2_signals[0][7][19] , 
        \s_mux2_signals[0][7][18] , \s_mux2_signals[0][7][17] , 
        \s_mux2_signals[0][7][16] , \s_mux2_signals[0][7][15] , 
        \s_mux2_signals[0][7][14] , \s_mux2_signals[0][7][13] , 
        \s_mux2_signals[0][7][12] , \s_mux2_signals[0][7][11] , 
        \s_mux2_signals[0][7][10] , \s_mux2_signals[0][7][9] , 
        \s_mux2_signals[0][7][8] , \s_mux2_signals[0][7][7] , 
        \s_mux2_signals[0][7][6] , \s_mux2_signals[0][7][5] , 
        \s_mux2_signals[0][7][4] , \s_mux2_signals[0][7][3] , 
        \s_mux2_signals[0][7][2] , \s_mux2_signals[0][7][1] , 
        \s_mux2_signals[0][7][0] }), .sel(n22), .portY({
        \s_mux1_signals[1][6][31] , \s_mux1_signals[1][6][30] , 
        \s_mux1_signals[1][6][29] , \s_mux1_signals[1][6][28] , 
        \s_mux1_signals[1][6][27] , \s_mux1_signals[1][6][26] , 
        \s_mux1_signals[1][6][25] , \s_mux1_signals[1][6][24] , 
        \s_mux1_signals[1][6][23] , \s_mux1_signals[1][6][22] , 
        \s_mux1_signals[1][6][21] , \s_mux1_signals[1][6][20] , 
        \s_mux1_signals[1][6][19] , \s_mux1_signals[1][6][18] , 
        \s_mux1_signals[1][6][17] , \s_mux1_signals[1][6][16] , 
        \s_mux1_signals[1][6][15] , \s_mux1_signals[1][6][14] , 
        \s_mux1_signals[1][6][13] , \s_mux1_signals[1][6][12] , 
        \s_mux1_signals[1][6][11] , \s_mux1_signals[1][6][10] , 
        \s_mux1_signals[1][6][9] , \s_mux1_signals[1][6][8] , 
        \s_mux1_signals[1][6][7] , \s_mux1_signals[1][6][6] , 
        \s_mux1_signals[1][6][5] , \s_mux1_signals[1][6][4] , 
        \s_mux1_signals[1][6][3] , \s_mux1_signals[1][6][2] , 
        \s_mux1_signals[1][6][1] , \s_mux1_signals[1][6][0] }) );
  Mux_NBit_2x1_NBIT_IN32_75 MUX1_0_8 ( .port0({\s_mux2_signals[0][8][31] , 
        \s_mux2_signals[0][8][30] , \s_mux2_signals[0][8][29] , 
        \s_mux2_signals[0][8][28] , \s_mux2_signals[0][8][27] , 
        \s_mux2_signals[0][8][26] , \s_mux2_signals[0][8][25] , 
        \s_mux2_signals[0][8][24] , \s_mux2_signals[0][8][23] , 
        \s_mux2_signals[0][8][22] , \s_mux2_signals[0][8][21] , 
        \s_mux2_signals[0][8][20] , \s_mux2_signals[0][8][19] , 
        \s_mux2_signals[0][8][18] , \s_mux2_signals[0][8][17] , 
        \s_mux2_signals[0][8][16] , \s_mux2_signals[0][8][15] , 
        \s_mux2_signals[0][8][14] , \s_mux2_signals[0][8][13] , 
        \s_mux2_signals[0][8][12] , \s_mux2_signals[0][8][11] , 
        \s_mux2_signals[0][8][10] , \s_mux2_signals[0][8][9] , 
        \s_mux2_signals[0][8][8] , \s_mux2_signals[0][8][7] , 
        \s_mux2_signals[0][8][6] , \s_mux2_signals[0][8][5] , 
        \s_mux2_signals[0][8][4] , \s_mux2_signals[0][8][3] , 
        \s_mux2_signals[0][8][2] , \s_mux2_signals[0][8][1] , 
        \s_mux2_signals[0][8][0] }), .port1({\s_mux2_signals[0][9][31] , 
        \s_mux2_signals[0][9][30] , \s_mux2_signals[0][9][29] , 
        \s_mux2_signals[0][9][28] , \s_mux2_signals[0][9][27] , 
        \s_mux2_signals[0][9][26] , \s_mux2_signals[0][9][25] , 
        \s_mux2_signals[0][9][24] , \s_mux2_signals[0][9][23] , 
        \s_mux2_signals[0][9][22] , \s_mux2_signals[0][9][21] , 
        \s_mux2_signals[0][9][20] , \s_mux2_signals[0][9][19] , 
        \s_mux2_signals[0][9][18] , \s_mux2_signals[0][9][17] , 
        \s_mux2_signals[0][9][16] , \s_mux2_signals[0][9][15] , 
        \s_mux2_signals[0][9][14] , \s_mux2_signals[0][9][13] , 
        \s_mux2_signals[0][9][12] , \s_mux2_signals[0][9][11] , 
        \s_mux2_signals[0][9][10] , \s_mux2_signals[0][9][9] , 
        \s_mux2_signals[0][9][8] , \s_mux2_signals[0][9][7] , 
        \s_mux2_signals[0][9][6] , \s_mux2_signals[0][9][5] , 
        \s_mux2_signals[0][9][4] , \s_mux2_signals[0][9][3] , 
        \s_mux2_signals[0][9][2] , \s_mux2_signals[0][9][1] , 
        \s_mux2_signals[0][9][0] }), .sel(n22), .portY({
        \s_mux1_signals[1][8][31] , \s_mux1_signals[1][8][30] , 
        \s_mux1_signals[1][8][29] , \s_mux1_signals[1][8][28] , 
        \s_mux1_signals[1][8][27] , \s_mux1_signals[1][8][26] , 
        \s_mux1_signals[1][8][25] , \s_mux1_signals[1][8][24] , 
        \s_mux1_signals[1][8][23] , \s_mux1_signals[1][8][22] , 
        \s_mux1_signals[1][8][21] , \s_mux1_signals[1][8][20] , 
        \s_mux1_signals[1][8][19] , \s_mux1_signals[1][8][18] , 
        \s_mux1_signals[1][8][17] , \s_mux1_signals[1][8][16] , 
        \s_mux1_signals[1][8][15] , \s_mux1_signals[1][8][14] , 
        \s_mux1_signals[1][8][13] , \s_mux1_signals[1][8][12] , 
        \s_mux1_signals[1][8][11] , \s_mux1_signals[1][8][10] , 
        \s_mux1_signals[1][8][9] , \s_mux1_signals[1][8][8] , 
        \s_mux1_signals[1][8][7] , \s_mux1_signals[1][8][6] , 
        \s_mux1_signals[1][8][5] , \s_mux1_signals[1][8][4] , 
        \s_mux1_signals[1][8][3] , \s_mux1_signals[1][8][2] , 
        \s_mux1_signals[1][8][1] , \s_mux1_signals[1][8][0] }) );
  Mux_NBit_2x1_NBIT_IN32_74 MUX1_0_10 ( .port0({\s_mux2_signals[0][10][31] , 
        \s_mux2_signals[0][10][30] , \s_mux2_signals[0][10][29] , 
        \s_mux2_signals[0][10][28] , \s_mux2_signals[0][10][27] , 
        \s_mux2_signals[0][10][26] , \s_mux2_signals[0][10][25] , 
        \s_mux2_signals[0][10][24] , \s_mux2_signals[0][10][23] , 
        \s_mux2_signals[0][10][22] , \s_mux2_signals[0][10][21] , 
        \s_mux2_signals[0][10][20] , \s_mux2_signals[0][10][19] , 
        \s_mux2_signals[0][10][18] , \s_mux2_signals[0][10][17] , 
        \s_mux2_signals[0][10][16] , \s_mux2_signals[0][10][15] , 
        \s_mux2_signals[0][10][14] , \s_mux2_signals[0][10][13] , 
        \s_mux2_signals[0][10][12] , \s_mux2_signals[0][10][11] , 
        \s_mux2_signals[0][10][10] , \s_mux2_signals[0][10][9] , 
        \s_mux2_signals[0][10][8] , \s_mux2_signals[0][10][7] , 
        \s_mux2_signals[0][10][6] , \s_mux2_signals[0][10][5] , 
        \s_mux2_signals[0][10][4] , \s_mux2_signals[0][10][3] , 
        \s_mux2_signals[0][10][2] , \s_mux2_signals[0][10][1] , 
        \s_mux2_signals[0][10][0] }), .port1({\s_mux2_signals[0][11][31] , 
        \s_mux2_signals[0][11][30] , \s_mux2_signals[0][11][29] , 
        \s_mux2_signals[0][11][28] , \s_mux2_signals[0][11][27] , 
        \s_mux2_signals[0][11][26] , \s_mux2_signals[0][11][25] , 
        \s_mux2_signals[0][11][24] , \s_mux2_signals[0][11][23] , 
        \s_mux2_signals[0][11][22] , \s_mux2_signals[0][11][21] , 
        \s_mux2_signals[0][11][20] , \s_mux2_signals[0][11][19] , 
        \s_mux2_signals[0][11][18] , \s_mux2_signals[0][11][17] , 
        \s_mux2_signals[0][11][16] , \s_mux2_signals[0][11][15] , 
        \s_mux2_signals[0][11][14] , \s_mux2_signals[0][11][13] , 
        \s_mux2_signals[0][11][12] , \s_mux2_signals[0][11][11] , 
        \s_mux2_signals[0][11][10] , \s_mux2_signals[0][11][9] , 
        \s_mux2_signals[0][11][8] , \s_mux2_signals[0][11][7] , 
        \s_mux2_signals[0][11][6] , \s_mux2_signals[0][11][5] , 
        \s_mux2_signals[0][11][4] , \s_mux2_signals[0][11][3] , 
        \s_mux2_signals[0][11][2] , \s_mux2_signals[0][11][1] , 
        \s_mux2_signals[0][11][0] }), .sel(n22), .portY({
        \s_mux1_signals[1][10][31] , \s_mux1_signals[1][10][30] , 
        \s_mux1_signals[1][10][29] , \s_mux1_signals[1][10][28] , 
        \s_mux1_signals[1][10][27] , \s_mux1_signals[1][10][26] , 
        \s_mux1_signals[1][10][25] , \s_mux1_signals[1][10][24] , 
        \s_mux1_signals[1][10][23] , \s_mux1_signals[1][10][22] , 
        \s_mux1_signals[1][10][21] , \s_mux1_signals[1][10][20] , 
        \s_mux1_signals[1][10][19] , \s_mux1_signals[1][10][18] , 
        \s_mux1_signals[1][10][17] , \s_mux1_signals[1][10][16] , 
        \s_mux1_signals[1][10][15] , \s_mux1_signals[1][10][14] , 
        \s_mux1_signals[1][10][13] , \s_mux1_signals[1][10][12] , 
        \s_mux1_signals[1][10][11] , \s_mux1_signals[1][10][10] , 
        \s_mux1_signals[1][10][9] , \s_mux1_signals[1][10][8] , 
        \s_mux1_signals[1][10][7] , \s_mux1_signals[1][10][6] , 
        \s_mux1_signals[1][10][5] , \s_mux1_signals[1][10][4] , 
        \s_mux1_signals[1][10][3] , \s_mux1_signals[1][10][2] , 
        \s_mux1_signals[1][10][1] , \s_mux1_signals[1][10][0] }) );
  Mux_NBit_2x1_NBIT_IN32_73 MUX1_0_12 ( .port0({\s_mux2_signals[0][12][31] , 
        \s_mux2_signals[0][12][30] , \s_mux2_signals[0][12][29] , 
        \s_mux2_signals[0][12][28] , \s_mux2_signals[0][12][27] , 
        \s_mux2_signals[0][12][26] , \s_mux2_signals[0][12][25] , 
        \s_mux2_signals[0][12][24] , \s_mux2_signals[0][12][23] , 
        \s_mux2_signals[0][12][22] , \s_mux2_signals[0][12][21] , 
        \s_mux2_signals[0][12][20] , \s_mux2_signals[0][12][19] , 
        \s_mux2_signals[0][12][18] , \s_mux2_signals[0][12][17] , 
        \s_mux2_signals[0][12][16] , \s_mux2_signals[0][12][15] , 
        \s_mux2_signals[0][12][14] , \s_mux2_signals[0][12][13] , 
        \s_mux2_signals[0][12][12] , \s_mux2_signals[0][12][11] , 
        \s_mux2_signals[0][12][10] , \s_mux2_signals[0][12][9] , 
        \s_mux2_signals[0][12][8] , \s_mux2_signals[0][12][7] , 
        \s_mux2_signals[0][12][6] , \s_mux2_signals[0][12][5] , 
        \s_mux2_signals[0][12][4] , \s_mux2_signals[0][12][3] , 
        \s_mux2_signals[0][12][2] , \s_mux2_signals[0][12][1] , 
        \s_mux2_signals[0][12][0] }), .port1({\s_mux2_signals[0][13][31] , 
        \s_mux2_signals[0][13][30] , \s_mux2_signals[0][13][29] , 
        \s_mux2_signals[0][13][28] , \s_mux2_signals[0][13][27] , 
        \s_mux2_signals[0][13][26] , \s_mux2_signals[0][13][25] , 
        \s_mux2_signals[0][13][24] , \s_mux2_signals[0][13][23] , 
        \s_mux2_signals[0][13][22] , \s_mux2_signals[0][13][21] , 
        \s_mux2_signals[0][13][20] , \s_mux2_signals[0][13][19] , 
        \s_mux2_signals[0][13][18] , \s_mux2_signals[0][13][17] , 
        \s_mux2_signals[0][13][16] , \s_mux2_signals[0][13][15] , 
        \s_mux2_signals[0][13][14] , \s_mux2_signals[0][13][13] , 
        \s_mux2_signals[0][13][12] , \s_mux2_signals[0][13][11] , 
        \s_mux2_signals[0][13][10] , \s_mux2_signals[0][13][9] , 
        \s_mux2_signals[0][13][8] , \s_mux2_signals[0][13][7] , 
        \s_mux2_signals[0][13][6] , \s_mux2_signals[0][13][5] , 
        \s_mux2_signals[0][13][4] , \s_mux2_signals[0][13][3] , 
        \s_mux2_signals[0][13][2] , \s_mux2_signals[0][13][1] , 
        \s_mux2_signals[0][13][0] }), .sel(n23), .portY({
        \s_mux1_signals[1][12][31] , \s_mux1_signals[1][12][30] , 
        \s_mux1_signals[1][12][29] , \s_mux1_signals[1][12][28] , 
        \s_mux1_signals[1][12][27] , \s_mux1_signals[1][12][26] , 
        \s_mux1_signals[1][12][25] , \s_mux1_signals[1][12][24] , 
        \s_mux1_signals[1][12][23] , \s_mux1_signals[1][12][22] , 
        \s_mux1_signals[1][12][21] , \s_mux1_signals[1][12][20] , 
        \s_mux1_signals[1][12][19] , \s_mux1_signals[1][12][18] , 
        \s_mux1_signals[1][12][17] , \s_mux1_signals[1][12][16] , 
        \s_mux1_signals[1][12][15] , \s_mux1_signals[1][12][14] , 
        \s_mux1_signals[1][12][13] , \s_mux1_signals[1][12][12] , 
        \s_mux1_signals[1][12][11] , \s_mux1_signals[1][12][10] , 
        \s_mux1_signals[1][12][9] , \s_mux1_signals[1][12][8] , 
        \s_mux1_signals[1][12][7] , \s_mux1_signals[1][12][6] , 
        \s_mux1_signals[1][12][5] , \s_mux1_signals[1][12][4] , 
        \s_mux1_signals[1][12][3] , \s_mux1_signals[1][12][2] , 
        \s_mux1_signals[1][12][1] , \s_mux1_signals[1][12][0] }) );
  Mux_NBit_2x1_NBIT_IN32_72 MUX1_0_14 ( .port0({\s_mux2_signals[0][14][31] , 
        \s_mux2_signals[0][14][30] , \s_mux2_signals[0][14][29] , 
        \s_mux2_signals[0][14][28] , \s_mux2_signals[0][14][27] , 
        \s_mux2_signals[0][14][26] , \s_mux2_signals[0][14][25] , 
        \s_mux2_signals[0][14][24] , \s_mux2_signals[0][14][23] , 
        \s_mux2_signals[0][14][22] , \s_mux2_signals[0][14][21] , 
        \s_mux2_signals[0][14][20] , \s_mux2_signals[0][14][19] , 
        \s_mux2_signals[0][14][18] , \s_mux2_signals[0][14][17] , 
        \s_mux2_signals[0][14][16] , \s_mux2_signals[0][14][15] , 
        \s_mux2_signals[0][14][14] , \s_mux2_signals[0][14][13] , 
        \s_mux2_signals[0][14][12] , \s_mux2_signals[0][14][11] , 
        \s_mux2_signals[0][14][10] , \s_mux2_signals[0][14][9] , 
        \s_mux2_signals[0][14][8] , \s_mux2_signals[0][14][7] , 
        \s_mux2_signals[0][14][6] , \s_mux2_signals[0][14][5] , 
        \s_mux2_signals[0][14][4] , \s_mux2_signals[0][14][3] , 
        \s_mux2_signals[0][14][2] , \s_mux2_signals[0][14][1] , 
        \s_mux2_signals[0][14][0] }), .port1({\s_mux2_signals[0][15][31] , 
        \s_mux2_signals[0][15][30] , \s_mux2_signals[0][15][29] , 
        \s_mux2_signals[0][15][28] , \s_mux2_signals[0][15][27] , 
        \s_mux2_signals[0][15][26] , \s_mux2_signals[0][15][25] , 
        \s_mux2_signals[0][15][24] , \s_mux2_signals[0][15][23] , 
        \s_mux2_signals[0][15][22] , \s_mux2_signals[0][15][21] , 
        \s_mux2_signals[0][15][20] , \s_mux2_signals[0][15][19] , 
        \s_mux2_signals[0][15][18] , \s_mux2_signals[0][15][17] , 
        \s_mux2_signals[0][15][16] , \s_mux2_signals[0][15][15] , 
        \s_mux2_signals[0][15][14] , \s_mux2_signals[0][15][13] , 
        \s_mux2_signals[0][15][12] , \s_mux2_signals[0][15][11] , 
        \s_mux2_signals[0][15][10] , \s_mux2_signals[0][15][9] , 
        \s_mux2_signals[0][15][8] , \s_mux2_signals[0][15][7] , 
        \s_mux2_signals[0][15][6] , \s_mux2_signals[0][15][5] , 
        \s_mux2_signals[0][15][4] , \s_mux2_signals[0][15][3] , 
        \s_mux2_signals[0][15][2] , \s_mux2_signals[0][15][1] , 
        \s_mux2_signals[0][15][0] }), .sel(n22), .portY({
        \s_mux1_signals[1][14][31] , \s_mux1_signals[1][14][30] , 
        \s_mux1_signals[1][14][29] , \s_mux1_signals[1][14][28] , 
        \s_mux1_signals[1][14][27] , \s_mux1_signals[1][14][26] , 
        \s_mux1_signals[1][14][25] , \s_mux1_signals[1][14][24] , 
        \s_mux1_signals[1][14][23] , \s_mux1_signals[1][14][22] , 
        \s_mux1_signals[1][14][21] , \s_mux1_signals[1][14][20] , 
        \s_mux1_signals[1][14][19] , \s_mux1_signals[1][14][18] , 
        \s_mux1_signals[1][14][17] , \s_mux1_signals[1][14][16] , 
        \s_mux1_signals[1][14][15] , \s_mux1_signals[1][14][14] , 
        \s_mux1_signals[1][14][13] , \s_mux1_signals[1][14][12] , 
        \s_mux1_signals[1][14][11] , \s_mux1_signals[1][14][10] , 
        \s_mux1_signals[1][14][9] , \s_mux1_signals[1][14][8] , 
        \s_mux1_signals[1][14][7] , \s_mux1_signals[1][14][6] , 
        \s_mux1_signals[1][14][5] , \s_mux1_signals[1][14][4] , 
        \s_mux1_signals[1][14][3] , \s_mux1_signals[1][14][2] , 
        \s_mux1_signals[1][14][1] , \s_mux1_signals[1][14][0] }) );
  Mux_NBit_2x1_NBIT_IN32_71 MUX1_0_16 ( .port0({\s_mux2_signals[0][16][31] , 
        \s_mux2_signals[0][16][30] , \s_mux2_signals[0][16][29] , 
        \s_mux2_signals[0][16][28] , \s_mux2_signals[0][16][27] , 
        \s_mux2_signals[0][16][26] , \s_mux2_signals[0][16][25] , 
        \s_mux2_signals[0][16][24] , \s_mux2_signals[0][16][23] , 
        \s_mux2_signals[0][16][22] , \s_mux2_signals[0][16][21] , 
        \s_mux2_signals[0][16][20] , \s_mux2_signals[0][16][19] , 
        \s_mux2_signals[0][16][18] , \s_mux2_signals[0][16][17] , 
        \s_mux2_signals[0][16][16] , \s_mux2_signals[0][16][15] , 
        \s_mux2_signals[0][16][14] , \s_mux2_signals[0][16][13] , 
        \s_mux2_signals[0][16][12] , \s_mux2_signals[0][16][11] , 
        \s_mux2_signals[0][16][10] , \s_mux2_signals[0][16][9] , 
        \s_mux2_signals[0][16][8] , \s_mux2_signals[0][16][7] , 
        \s_mux2_signals[0][16][6] , \s_mux2_signals[0][16][5] , 
        \s_mux2_signals[0][16][4] , \s_mux2_signals[0][16][3] , 
        \s_mux2_signals[0][16][2] , \s_mux2_signals[0][16][1] , 
        \s_mux2_signals[0][16][0] }), .port1({\s_mux2_signals[0][17][31] , 
        \s_mux2_signals[0][17][30] , \s_mux2_signals[0][17][29] , 
        \s_mux2_signals[0][17][28] , \s_mux2_signals[0][17][27] , 
        \s_mux2_signals[0][17][26] , \s_mux2_signals[0][17][25] , 
        \s_mux2_signals[0][17][24] , \s_mux2_signals[0][17][23] , 
        \s_mux2_signals[0][17][22] , \s_mux2_signals[0][17][21] , 
        \s_mux2_signals[0][17][20] , \s_mux2_signals[0][17][19] , 
        \s_mux2_signals[0][17][18] , \s_mux2_signals[0][17][17] , 
        \s_mux2_signals[0][17][16] , \s_mux2_signals[0][17][15] , 
        \s_mux2_signals[0][17][14] , \s_mux2_signals[0][17][13] , 
        \s_mux2_signals[0][17][12] , \s_mux2_signals[0][17][11] , 
        \s_mux2_signals[0][17][10] , \s_mux2_signals[0][17][9] , 
        \s_mux2_signals[0][17][8] , \s_mux2_signals[0][17][7] , 
        \s_mux2_signals[0][17][6] , \s_mux2_signals[0][17][5] , 
        \s_mux2_signals[0][17][4] , \s_mux2_signals[0][17][3] , 
        \s_mux2_signals[0][17][2] , \s_mux2_signals[0][17][1] , 
        \s_mux2_signals[0][17][0] }), .sel(n23), .portY({
        \s_mux1_signals[1][16][31] , \s_mux1_signals[1][16][30] , 
        \s_mux1_signals[1][16][29] , \s_mux1_signals[1][16][28] , 
        \s_mux1_signals[1][16][27] , \s_mux1_signals[1][16][26] , 
        \s_mux1_signals[1][16][25] , \s_mux1_signals[1][16][24] , 
        \s_mux1_signals[1][16][23] , \s_mux1_signals[1][16][22] , 
        \s_mux1_signals[1][16][21] , \s_mux1_signals[1][16][20] , 
        \s_mux1_signals[1][16][19] , \s_mux1_signals[1][16][18] , 
        \s_mux1_signals[1][16][17] , \s_mux1_signals[1][16][16] , 
        \s_mux1_signals[1][16][15] , \s_mux1_signals[1][16][14] , 
        \s_mux1_signals[1][16][13] , \s_mux1_signals[1][16][12] , 
        \s_mux1_signals[1][16][11] , \s_mux1_signals[1][16][10] , 
        \s_mux1_signals[1][16][9] , \s_mux1_signals[1][16][8] , 
        \s_mux1_signals[1][16][7] , \s_mux1_signals[1][16][6] , 
        \s_mux1_signals[1][16][5] , \s_mux1_signals[1][16][4] , 
        \s_mux1_signals[1][16][3] , \s_mux1_signals[1][16][2] , 
        \s_mux1_signals[1][16][1] , \s_mux1_signals[1][16][0] }) );
  Mux_NBit_2x1_NBIT_IN32_70 MUX1_0_18 ( .port0({\s_mux2_signals[0][18][31] , 
        \s_mux2_signals[0][18][30] , \s_mux2_signals[0][18][29] , 
        \s_mux2_signals[0][18][28] , \s_mux2_signals[0][18][27] , 
        \s_mux2_signals[0][18][26] , \s_mux2_signals[0][18][25] , 
        \s_mux2_signals[0][18][24] , \s_mux2_signals[0][18][23] , 
        \s_mux2_signals[0][18][22] , \s_mux2_signals[0][18][21] , 
        \s_mux2_signals[0][18][20] , \s_mux2_signals[0][18][19] , 
        \s_mux2_signals[0][18][18] , \s_mux2_signals[0][18][17] , 
        \s_mux2_signals[0][18][16] , \s_mux2_signals[0][18][15] , 
        \s_mux2_signals[0][18][14] , \s_mux2_signals[0][18][13] , 
        \s_mux2_signals[0][18][12] , \s_mux2_signals[0][18][11] , 
        \s_mux2_signals[0][18][10] , \s_mux2_signals[0][18][9] , 
        \s_mux2_signals[0][18][8] , \s_mux2_signals[0][18][7] , 
        \s_mux2_signals[0][18][6] , \s_mux2_signals[0][18][5] , 
        \s_mux2_signals[0][18][4] , \s_mux2_signals[0][18][3] , 
        \s_mux2_signals[0][18][2] , \s_mux2_signals[0][18][1] , 
        \s_mux2_signals[0][18][0] }), .port1({\s_mux2_signals[0][19][31] , 
        \s_mux2_signals[0][19][30] , \s_mux2_signals[0][19][29] , 
        \s_mux2_signals[0][19][28] , \s_mux2_signals[0][19][27] , 
        \s_mux2_signals[0][19][26] , \s_mux2_signals[0][19][25] , 
        \s_mux2_signals[0][19][24] , \s_mux2_signals[0][19][23] , 
        \s_mux2_signals[0][19][22] , \s_mux2_signals[0][19][21] , 
        \s_mux2_signals[0][19][20] , \s_mux2_signals[0][19][19] , 
        \s_mux2_signals[0][19][18] , \s_mux2_signals[0][19][17] , 
        \s_mux2_signals[0][19][16] , \s_mux2_signals[0][19][15] , 
        \s_mux2_signals[0][19][14] , \s_mux2_signals[0][19][13] , 
        \s_mux2_signals[0][19][12] , \s_mux2_signals[0][19][11] , 
        \s_mux2_signals[0][19][10] , \s_mux2_signals[0][19][9] , 
        \s_mux2_signals[0][19][8] , \s_mux2_signals[0][19][7] , 
        \s_mux2_signals[0][19][6] , \s_mux2_signals[0][19][5] , 
        \s_mux2_signals[0][19][4] , \s_mux2_signals[0][19][3] , 
        \s_mux2_signals[0][19][2] , \s_mux2_signals[0][19][1] , 
        \s_mux2_signals[0][19][0] }), .sel(n23), .portY({
        \s_mux1_signals[1][18][31] , \s_mux1_signals[1][18][30] , 
        \s_mux1_signals[1][18][29] , \s_mux1_signals[1][18][28] , 
        \s_mux1_signals[1][18][27] , \s_mux1_signals[1][18][26] , 
        \s_mux1_signals[1][18][25] , \s_mux1_signals[1][18][24] , 
        \s_mux1_signals[1][18][23] , \s_mux1_signals[1][18][22] , 
        \s_mux1_signals[1][18][21] , \s_mux1_signals[1][18][20] , 
        \s_mux1_signals[1][18][19] , \s_mux1_signals[1][18][18] , 
        \s_mux1_signals[1][18][17] , \s_mux1_signals[1][18][16] , 
        \s_mux1_signals[1][18][15] , \s_mux1_signals[1][18][14] , 
        \s_mux1_signals[1][18][13] , \s_mux1_signals[1][18][12] , 
        \s_mux1_signals[1][18][11] , \s_mux1_signals[1][18][10] , 
        \s_mux1_signals[1][18][9] , \s_mux1_signals[1][18][8] , 
        \s_mux1_signals[1][18][7] , \s_mux1_signals[1][18][6] , 
        \s_mux1_signals[1][18][5] , \s_mux1_signals[1][18][4] , 
        \s_mux1_signals[1][18][3] , \s_mux1_signals[1][18][2] , 
        \s_mux1_signals[1][18][1] , \s_mux1_signals[1][18][0] }) );
  Mux_NBit_2x1_NBIT_IN32_69 MUX1_0_20 ( .port0({\s_mux2_signals[0][20][31] , 
        \s_mux2_signals[0][20][30] , \s_mux2_signals[0][20][29] , 
        \s_mux2_signals[0][20][28] , \s_mux2_signals[0][20][27] , 
        \s_mux2_signals[0][20][26] , \s_mux2_signals[0][20][25] , 
        \s_mux2_signals[0][20][24] , \s_mux2_signals[0][20][23] , 
        \s_mux2_signals[0][20][22] , \s_mux2_signals[0][20][21] , 
        \s_mux2_signals[0][20][20] , \s_mux2_signals[0][20][19] , 
        \s_mux2_signals[0][20][18] , \s_mux2_signals[0][20][17] , 
        \s_mux2_signals[0][20][16] , \s_mux2_signals[0][20][15] , 
        \s_mux2_signals[0][20][14] , \s_mux2_signals[0][20][13] , 
        \s_mux2_signals[0][20][12] , \s_mux2_signals[0][20][11] , 
        \s_mux2_signals[0][20][10] , \s_mux2_signals[0][20][9] , 
        \s_mux2_signals[0][20][8] , \s_mux2_signals[0][20][7] , 
        \s_mux2_signals[0][20][6] , \s_mux2_signals[0][20][5] , 
        \s_mux2_signals[0][20][4] , \s_mux2_signals[0][20][3] , 
        \s_mux2_signals[0][20][2] , \s_mux2_signals[0][20][1] , 
        \s_mux2_signals[0][20][0] }), .port1({\s_mux2_signals[0][21][31] , 
        \s_mux2_signals[0][21][30] , \s_mux2_signals[0][21][29] , 
        \s_mux2_signals[0][21][28] , \s_mux2_signals[0][21][27] , 
        \s_mux2_signals[0][21][26] , \s_mux2_signals[0][21][25] , 
        \s_mux2_signals[0][21][24] , \s_mux2_signals[0][21][23] , 
        \s_mux2_signals[0][21][22] , \s_mux2_signals[0][21][21] , 
        \s_mux2_signals[0][21][20] , \s_mux2_signals[0][21][19] , 
        \s_mux2_signals[0][21][18] , \s_mux2_signals[0][21][17] , 
        \s_mux2_signals[0][21][16] , \s_mux2_signals[0][21][15] , 
        \s_mux2_signals[0][21][14] , \s_mux2_signals[0][21][13] , 
        \s_mux2_signals[0][21][12] , \s_mux2_signals[0][21][11] , 
        \s_mux2_signals[0][21][10] , \s_mux2_signals[0][21][9] , 
        \s_mux2_signals[0][21][8] , \s_mux2_signals[0][21][7] , 
        \s_mux2_signals[0][21][6] , \s_mux2_signals[0][21][5] , 
        \s_mux2_signals[0][21][4] , \s_mux2_signals[0][21][3] , 
        \s_mux2_signals[0][21][2] , \s_mux2_signals[0][21][1] , 
        \s_mux2_signals[0][21][0] }), .sel(n23), .portY({
        \s_mux1_signals[1][20][31] , \s_mux1_signals[1][20][30] , 
        \s_mux1_signals[1][20][29] , \s_mux1_signals[1][20][28] , 
        \s_mux1_signals[1][20][27] , \s_mux1_signals[1][20][26] , 
        \s_mux1_signals[1][20][25] , \s_mux1_signals[1][20][24] , 
        \s_mux1_signals[1][20][23] , \s_mux1_signals[1][20][22] , 
        \s_mux1_signals[1][20][21] , \s_mux1_signals[1][20][20] , 
        \s_mux1_signals[1][20][19] , \s_mux1_signals[1][20][18] , 
        \s_mux1_signals[1][20][17] , \s_mux1_signals[1][20][16] , 
        \s_mux1_signals[1][20][15] , \s_mux1_signals[1][20][14] , 
        \s_mux1_signals[1][20][13] , \s_mux1_signals[1][20][12] , 
        \s_mux1_signals[1][20][11] , \s_mux1_signals[1][20][10] , 
        \s_mux1_signals[1][20][9] , \s_mux1_signals[1][20][8] , 
        \s_mux1_signals[1][20][7] , \s_mux1_signals[1][20][6] , 
        \s_mux1_signals[1][20][5] , \s_mux1_signals[1][20][4] , 
        \s_mux1_signals[1][20][3] , \s_mux1_signals[1][20][2] , 
        \s_mux1_signals[1][20][1] , \s_mux1_signals[1][20][0] }) );
  Mux_NBit_2x1_NBIT_IN32_68 MUX1_0_22 ( .port0({\s_mux2_signals[0][22][31] , 
        \s_mux2_signals[0][22][30] , \s_mux2_signals[0][22][29] , 
        \s_mux2_signals[0][22][28] , \s_mux2_signals[0][22][27] , 
        \s_mux2_signals[0][22][26] , \s_mux2_signals[0][22][25] , 
        \s_mux2_signals[0][22][24] , \s_mux2_signals[0][22][23] , 
        \s_mux2_signals[0][22][22] , \s_mux2_signals[0][22][21] , 
        \s_mux2_signals[0][22][20] , \s_mux2_signals[0][22][19] , 
        \s_mux2_signals[0][22][18] , \s_mux2_signals[0][22][17] , 
        \s_mux2_signals[0][22][16] , \s_mux2_signals[0][22][15] , 
        \s_mux2_signals[0][22][14] , \s_mux2_signals[0][22][13] , 
        \s_mux2_signals[0][22][12] , \s_mux2_signals[0][22][11] , 
        \s_mux2_signals[0][22][10] , \s_mux2_signals[0][22][9] , 
        \s_mux2_signals[0][22][8] , \s_mux2_signals[0][22][7] , 
        \s_mux2_signals[0][22][6] , \s_mux2_signals[0][22][5] , 
        \s_mux2_signals[0][22][4] , \s_mux2_signals[0][22][3] , 
        \s_mux2_signals[0][22][2] , \s_mux2_signals[0][22][1] , 
        \s_mux2_signals[0][22][0] }), .port1({\s_mux2_signals[0][23][31] , 
        \s_mux2_signals[0][23][30] , \s_mux2_signals[0][23][29] , 
        \s_mux2_signals[0][23][28] , \s_mux2_signals[0][23][27] , 
        \s_mux2_signals[0][23][26] , \s_mux2_signals[0][23][25] , 
        \s_mux2_signals[0][23][24] , \s_mux2_signals[0][23][23] , 
        \s_mux2_signals[0][23][22] , \s_mux2_signals[0][23][21] , 
        \s_mux2_signals[0][23][20] , \s_mux2_signals[0][23][19] , 
        \s_mux2_signals[0][23][18] , \s_mux2_signals[0][23][17] , 
        \s_mux2_signals[0][23][16] , \s_mux2_signals[0][23][15] , 
        \s_mux2_signals[0][23][14] , \s_mux2_signals[0][23][13] , 
        \s_mux2_signals[0][23][12] , \s_mux2_signals[0][23][11] , 
        \s_mux2_signals[0][23][10] , \s_mux2_signals[0][23][9] , 
        \s_mux2_signals[0][23][8] , \s_mux2_signals[0][23][7] , 
        \s_mux2_signals[0][23][6] , \s_mux2_signals[0][23][5] , 
        \s_mux2_signals[0][23][4] , \s_mux2_signals[0][23][3] , 
        \s_mux2_signals[0][23][2] , \s_mux2_signals[0][23][1] , 
        \s_mux2_signals[0][23][0] }), .sel(n22), .portY({
        \s_mux1_signals[1][22][31] , \s_mux1_signals[1][22][30] , 
        \s_mux1_signals[1][22][29] , \s_mux1_signals[1][22][28] , 
        \s_mux1_signals[1][22][27] , \s_mux1_signals[1][22][26] , 
        \s_mux1_signals[1][22][25] , \s_mux1_signals[1][22][24] , 
        \s_mux1_signals[1][22][23] , \s_mux1_signals[1][22][22] , 
        \s_mux1_signals[1][22][21] , \s_mux1_signals[1][22][20] , 
        \s_mux1_signals[1][22][19] , \s_mux1_signals[1][22][18] , 
        \s_mux1_signals[1][22][17] , \s_mux1_signals[1][22][16] , 
        \s_mux1_signals[1][22][15] , \s_mux1_signals[1][22][14] , 
        \s_mux1_signals[1][22][13] , \s_mux1_signals[1][22][12] , 
        \s_mux1_signals[1][22][11] , \s_mux1_signals[1][22][10] , 
        \s_mux1_signals[1][22][9] , \s_mux1_signals[1][22][8] , 
        \s_mux1_signals[1][22][7] , \s_mux1_signals[1][22][6] , 
        \s_mux1_signals[1][22][5] , \s_mux1_signals[1][22][4] , 
        \s_mux1_signals[1][22][3] , \s_mux1_signals[1][22][2] , 
        \s_mux1_signals[1][22][1] , \s_mux1_signals[1][22][0] }) );
  Mux_NBit_2x1_NBIT_IN32_67 MUX1_0_24 ( .port0({\s_mux2_signals[0][24][31] , 
        \s_mux2_signals[0][24][30] , \s_mux2_signals[0][24][29] , 
        \s_mux2_signals[0][24][28] , \s_mux2_signals[0][24][27] , 
        \s_mux2_signals[0][24][26] , \s_mux2_signals[0][24][25] , 
        \s_mux2_signals[0][24][24] , \s_mux2_signals[0][24][23] , 
        \s_mux2_signals[0][24][22] , \s_mux2_signals[0][24][21] , 
        \s_mux2_signals[0][24][20] , \s_mux2_signals[0][24][19] , 
        \s_mux2_signals[0][24][18] , \s_mux2_signals[0][24][17] , 
        \s_mux2_signals[0][24][16] , \s_mux2_signals[0][24][15] , 
        \s_mux2_signals[0][24][14] , \s_mux2_signals[0][24][13] , 
        \s_mux2_signals[0][24][12] , \s_mux2_signals[0][24][11] , 
        \s_mux2_signals[0][24][10] , \s_mux2_signals[0][24][9] , 
        \s_mux2_signals[0][24][8] , \s_mux2_signals[0][24][7] , 
        \s_mux2_signals[0][24][6] , \s_mux2_signals[0][24][5] , 
        \s_mux2_signals[0][24][4] , \s_mux2_signals[0][24][3] , 
        \s_mux2_signals[0][24][2] , \s_mux2_signals[0][24][1] , 
        \s_mux2_signals[0][24][0] }), .port1({\s_mux2_signals[0][25][31] , 
        \s_mux2_signals[0][25][30] , \s_mux2_signals[0][25][29] , 
        \s_mux2_signals[0][25][28] , \s_mux2_signals[0][25][27] , 
        \s_mux2_signals[0][25][26] , \s_mux2_signals[0][25][25] , 
        \s_mux2_signals[0][25][24] , \s_mux2_signals[0][25][23] , 
        \s_mux2_signals[0][25][22] , \s_mux2_signals[0][25][21] , 
        \s_mux2_signals[0][25][20] , \s_mux2_signals[0][25][19] , 
        \s_mux2_signals[0][25][18] , \s_mux2_signals[0][25][17] , 
        \s_mux2_signals[0][25][16] , \s_mux2_signals[0][25][15] , 
        \s_mux2_signals[0][25][14] , \s_mux2_signals[0][25][13] , 
        \s_mux2_signals[0][25][12] , \s_mux2_signals[0][25][11] , 
        \s_mux2_signals[0][25][10] , \s_mux2_signals[0][25][9] , 
        \s_mux2_signals[0][25][8] , \s_mux2_signals[0][25][7] , 
        \s_mux2_signals[0][25][6] , \s_mux2_signals[0][25][5] , 
        \s_mux2_signals[0][25][4] , \s_mux2_signals[0][25][3] , 
        \s_mux2_signals[0][25][2] , \s_mux2_signals[0][25][1] , 
        \s_mux2_signals[0][25][0] }), .sel(n23), .portY({
        \s_mux1_signals[1][24][31] , \s_mux1_signals[1][24][30] , 
        \s_mux1_signals[1][24][29] , \s_mux1_signals[1][24][28] , 
        \s_mux1_signals[1][24][27] , \s_mux1_signals[1][24][26] , 
        \s_mux1_signals[1][24][25] , \s_mux1_signals[1][24][24] , 
        \s_mux1_signals[1][24][23] , \s_mux1_signals[1][24][22] , 
        \s_mux1_signals[1][24][21] , \s_mux1_signals[1][24][20] , 
        \s_mux1_signals[1][24][19] , \s_mux1_signals[1][24][18] , 
        \s_mux1_signals[1][24][17] , \s_mux1_signals[1][24][16] , 
        \s_mux1_signals[1][24][15] , \s_mux1_signals[1][24][14] , 
        \s_mux1_signals[1][24][13] , \s_mux1_signals[1][24][12] , 
        \s_mux1_signals[1][24][11] , \s_mux1_signals[1][24][10] , 
        \s_mux1_signals[1][24][9] , \s_mux1_signals[1][24][8] , 
        \s_mux1_signals[1][24][7] , \s_mux1_signals[1][24][6] , 
        \s_mux1_signals[1][24][5] , \s_mux1_signals[1][24][4] , 
        \s_mux1_signals[1][24][3] , \s_mux1_signals[1][24][2] , 
        \s_mux1_signals[1][24][1] , \s_mux1_signals[1][24][0] }) );
  Mux_NBit_2x1_NBIT_IN32_66 MUX1_0_26 ( .port0({\s_mux2_signals[0][26][31] , 
        \s_mux2_signals[0][26][30] , \s_mux2_signals[0][26][29] , 
        \s_mux2_signals[0][26][28] , \s_mux2_signals[0][26][27] , 
        \s_mux2_signals[0][26][26] , \s_mux2_signals[0][26][25] , 
        \s_mux2_signals[0][26][24] , \s_mux2_signals[0][26][23] , 
        \s_mux2_signals[0][26][22] , \s_mux2_signals[0][26][21] , 
        \s_mux2_signals[0][26][20] , \s_mux2_signals[0][26][19] , 
        \s_mux2_signals[0][26][18] , \s_mux2_signals[0][26][17] , 
        \s_mux2_signals[0][26][16] , \s_mux2_signals[0][26][15] , 
        \s_mux2_signals[0][26][14] , \s_mux2_signals[0][26][13] , 
        \s_mux2_signals[0][26][12] , \s_mux2_signals[0][26][11] , 
        \s_mux2_signals[0][26][10] , \s_mux2_signals[0][26][9] , 
        \s_mux2_signals[0][26][8] , \s_mux2_signals[0][26][7] , 
        \s_mux2_signals[0][26][6] , \s_mux2_signals[0][26][5] , 
        \s_mux2_signals[0][26][4] , \s_mux2_signals[0][26][3] , 
        \s_mux2_signals[0][26][2] , \s_mux2_signals[0][26][1] , 
        \s_mux2_signals[0][26][0] }), .port1({\s_mux2_signals[0][27][31] , 
        \s_mux2_signals[0][27][30] , \s_mux2_signals[0][27][29] , 
        \s_mux2_signals[0][27][28] , \s_mux2_signals[0][27][27] , 
        \s_mux2_signals[0][27][26] , \s_mux2_signals[0][27][25] , 
        \s_mux2_signals[0][27][24] , \s_mux2_signals[0][27][23] , 
        \s_mux2_signals[0][27][22] , \s_mux2_signals[0][27][21] , 
        \s_mux2_signals[0][27][20] , \s_mux2_signals[0][27][19] , 
        \s_mux2_signals[0][27][18] , \s_mux2_signals[0][27][17] , 
        \s_mux2_signals[0][27][16] , \s_mux2_signals[0][27][15] , 
        \s_mux2_signals[0][27][14] , \s_mux2_signals[0][27][13] , 
        \s_mux2_signals[0][27][12] , \s_mux2_signals[0][27][11] , 
        \s_mux2_signals[0][27][10] , \s_mux2_signals[0][27][9] , 
        \s_mux2_signals[0][27][8] , \s_mux2_signals[0][27][7] , 
        \s_mux2_signals[0][27][6] , \s_mux2_signals[0][27][5] , 
        \s_mux2_signals[0][27][4] , \s_mux2_signals[0][27][3] , 
        \s_mux2_signals[0][27][2] , \s_mux2_signals[0][27][1] , 
        \s_mux2_signals[0][27][0] }), .sel(n23), .portY({
        \s_mux1_signals[1][26][31] , \s_mux1_signals[1][26][30] , 
        \s_mux1_signals[1][26][29] , \s_mux1_signals[1][26][28] , 
        \s_mux1_signals[1][26][27] , \s_mux1_signals[1][26][26] , 
        \s_mux1_signals[1][26][25] , \s_mux1_signals[1][26][24] , 
        \s_mux1_signals[1][26][23] , \s_mux1_signals[1][26][22] , 
        \s_mux1_signals[1][26][21] , \s_mux1_signals[1][26][20] , 
        \s_mux1_signals[1][26][19] , \s_mux1_signals[1][26][18] , 
        \s_mux1_signals[1][26][17] , \s_mux1_signals[1][26][16] , 
        \s_mux1_signals[1][26][15] , \s_mux1_signals[1][26][14] , 
        \s_mux1_signals[1][26][13] , \s_mux1_signals[1][26][12] , 
        \s_mux1_signals[1][26][11] , \s_mux1_signals[1][26][10] , 
        \s_mux1_signals[1][26][9] , \s_mux1_signals[1][26][8] , 
        \s_mux1_signals[1][26][7] , \s_mux1_signals[1][26][6] , 
        \s_mux1_signals[1][26][5] , \s_mux1_signals[1][26][4] , 
        \s_mux1_signals[1][26][3] , \s_mux1_signals[1][26][2] , 
        \s_mux1_signals[1][26][1] , \s_mux1_signals[1][26][0] }) );
  Mux_NBit_2x1_NBIT_IN32_65 MUX1_0_28 ( .port0({\s_mux2_signals[0][28][31] , 
        \s_mux2_signals[0][28][30] , \s_mux2_signals[0][28][29] , 
        \s_mux2_signals[0][28][28] , \s_mux2_signals[0][28][27] , 
        \s_mux2_signals[0][28][26] , \s_mux2_signals[0][28][25] , 
        \s_mux2_signals[0][28][24] , \s_mux2_signals[0][28][23] , 
        \s_mux2_signals[0][28][22] , \s_mux2_signals[0][28][21] , 
        \s_mux2_signals[0][28][20] , \s_mux2_signals[0][28][19] , 
        \s_mux2_signals[0][28][18] , \s_mux2_signals[0][28][17] , 
        \s_mux2_signals[0][28][16] , \s_mux2_signals[0][28][15] , 
        \s_mux2_signals[0][28][14] , \s_mux2_signals[0][28][13] , 
        \s_mux2_signals[0][28][12] , \s_mux2_signals[0][28][11] , 
        \s_mux2_signals[0][28][10] , \s_mux2_signals[0][28][9] , 
        \s_mux2_signals[0][28][8] , \s_mux2_signals[0][28][7] , 
        \s_mux2_signals[0][28][6] , \s_mux2_signals[0][28][5] , 
        \s_mux2_signals[0][28][4] , \s_mux2_signals[0][28][3] , 
        \s_mux2_signals[0][28][2] , \s_mux2_signals[0][28][1] , 
        \s_mux2_signals[0][28][0] }), .port1({\s_mux2_signals[0][29][31] , 
        \s_mux2_signals[0][29][30] , \s_mux2_signals[0][29][29] , 
        \s_mux2_signals[0][29][28] , \s_mux2_signals[0][29][27] , 
        \s_mux2_signals[0][29][26] , \s_mux2_signals[0][29][25] , 
        \s_mux2_signals[0][29][24] , \s_mux2_signals[0][29][23] , 
        \s_mux2_signals[0][29][22] , \s_mux2_signals[0][29][21] , 
        \s_mux2_signals[0][29][20] , \s_mux2_signals[0][29][19] , 
        \s_mux2_signals[0][29][18] , \s_mux2_signals[0][29][17] , 
        \s_mux2_signals[0][29][16] , \s_mux2_signals[0][29][15] , 
        \s_mux2_signals[0][29][14] , \s_mux2_signals[0][29][13] , 
        \s_mux2_signals[0][29][12] , \s_mux2_signals[0][29][11] , 
        \s_mux2_signals[0][29][10] , \s_mux2_signals[0][29][9] , 
        \s_mux2_signals[0][29][8] , \s_mux2_signals[0][29][7] , 
        \s_mux2_signals[0][29][6] , \s_mux2_signals[0][29][5] , 
        \s_mux2_signals[0][29][4] , \s_mux2_signals[0][29][3] , 
        \s_mux2_signals[0][29][2] , \s_mux2_signals[0][29][1] , 
        \s_mux2_signals[0][29][0] }), .sel(n23), .portY({
        \s_mux1_signals[1][28][31] , \s_mux1_signals[1][28][30] , 
        \s_mux1_signals[1][28][29] , \s_mux1_signals[1][28][28] , 
        \s_mux1_signals[1][28][27] , \s_mux1_signals[1][28][26] , 
        \s_mux1_signals[1][28][25] , \s_mux1_signals[1][28][24] , 
        \s_mux1_signals[1][28][23] , \s_mux1_signals[1][28][22] , 
        \s_mux1_signals[1][28][21] , \s_mux1_signals[1][28][20] , 
        \s_mux1_signals[1][28][19] , \s_mux1_signals[1][28][18] , 
        \s_mux1_signals[1][28][17] , \s_mux1_signals[1][28][16] , 
        \s_mux1_signals[1][28][15] , \s_mux1_signals[1][28][14] , 
        \s_mux1_signals[1][28][13] , \s_mux1_signals[1][28][12] , 
        \s_mux1_signals[1][28][11] , \s_mux1_signals[1][28][10] , 
        \s_mux1_signals[1][28][9] , \s_mux1_signals[1][28][8] , 
        \s_mux1_signals[1][28][7] , \s_mux1_signals[1][28][6] , 
        \s_mux1_signals[1][28][5] , \s_mux1_signals[1][28][4] , 
        \s_mux1_signals[1][28][3] , \s_mux1_signals[1][28][2] , 
        \s_mux1_signals[1][28][1] , \s_mux1_signals[1][28][0] }) );
  Mux_NBit_2x1_NBIT_IN32_64 MUX1_0_30 ( .port0({\s_mux2_signals[0][30][31] , 
        \s_mux2_signals[0][30][30] , \s_mux2_signals[0][30][29] , 
        \s_mux2_signals[0][30][28] , \s_mux2_signals[0][30][27] , 
        \s_mux2_signals[0][30][26] , \s_mux2_signals[0][30][25] , 
        \s_mux2_signals[0][30][24] , \s_mux2_signals[0][30][23] , 
        \s_mux2_signals[0][30][22] , \s_mux2_signals[0][30][21] , 
        \s_mux2_signals[0][30][20] , \s_mux2_signals[0][30][19] , 
        \s_mux2_signals[0][30][18] , \s_mux2_signals[0][30][17] , 
        \s_mux2_signals[0][30][16] , \s_mux2_signals[0][30][15] , 
        \s_mux2_signals[0][30][14] , \s_mux2_signals[0][30][13] , 
        \s_mux2_signals[0][30][12] , \s_mux2_signals[0][30][11] , 
        \s_mux2_signals[0][30][10] , \s_mux2_signals[0][30][9] , 
        \s_mux2_signals[0][30][8] , \s_mux2_signals[0][30][7] , 
        \s_mux2_signals[0][30][6] , \s_mux2_signals[0][30][5] , 
        \s_mux2_signals[0][30][4] , \s_mux2_signals[0][30][3] , 
        \s_mux2_signals[0][30][2] , \s_mux2_signals[0][30][1] , 
        \s_mux2_signals[0][30][0] }), .port1({\s_mux2_signals[0][31][31] , 
        \s_mux2_signals[0][31][30] , \s_mux2_signals[0][31][29] , 
        \s_mux2_signals[0][31][28] , \s_mux2_signals[0][31][27] , 
        \s_mux2_signals[0][31][26] , \s_mux2_signals[0][31][25] , 
        \s_mux2_signals[0][31][24] , \s_mux2_signals[0][31][23] , 
        \s_mux2_signals[0][31][22] , \s_mux2_signals[0][31][21] , 
        \s_mux2_signals[0][31][20] , \s_mux2_signals[0][31][19] , 
        \s_mux2_signals[0][31][18] , \s_mux2_signals[0][31][17] , 
        \s_mux2_signals[0][31][16] , \s_mux2_signals[0][31][15] , 
        \s_mux2_signals[0][31][14] , \s_mux2_signals[0][31][13] , 
        \s_mux2_signals[0][31][12] , \s_mux2_signals[0][31][11] , 
        \s_mux2_signals[0][31][10] , \s_mux2_signals[0][31][9] , 
        \s_mux2_signals[0][31][8] , \s_mux2_signals[0][31][7] , 
        \s_mux2_signals[0][31][6] , \s_mux2_signals[0][31][5] , 
        \s_mux2_signals[0][31][4] , \s_mux2_signals[0][31][3] , 
        \s_mux2_signals[0][31][2] , \s_mux2_signals[0][31][1] , 
        \s_mux2_signals[0][31][0] }), .sel(n24), .portY({
        \s_mux1_signals[1][30][31] , \s_mux1_signals[1][30][30] , 
        \s_mux1_signals[1][30][29] , \s_mux1_signals[1][30][28] , 
        \s_mux1_signals[1][30][27] , \s_mux1_signals[1][30][26] , 
        \s_mux1_signals[1][30][25] , \s_mux1_signals[1][30][24] , 
        \s_mux1_signals[1][30][23] , \s_mux1_signals[1][30][22] , 
        \s_mux1_signals[1][30][21] , \s_mux1_signals[1][30][20] , 
        \s_mux1_signals[1][30][19] , \s_mux1_signals[1][30][18] , 
        \s_mux1_signals[1][30][17] , \s_mux1_signals[1][30][16] , 
        \s_mux1_signals[1][30][15] , \s_mux1_signals[1][30][14] , 
        \s_mux1_signals[1][30][13] , \s_mux1_signals[1][30][12] , 
        \s_mux1_signals[1][30][11] , \s_mux1_signals[1][30][10] , 
        \s_mux1_signals[1][30][9] , \s_mux1_signals[1][30][8] , 
        \s_mux1_signals[1][30][7] , \s_mux1_signals[1][30][6] , 
        \s_mux1_signals[1][30][5] , \s_mux1_signals[1][30][4] , 
        \s_mux1_signals[1][30][3] , \s_mux1_signals[1][30][2] , 
        \s_mux1_signals[1][30][1] , \s_mux1_signals[1][30][0] }) );
  Mux_NBit_2x1_NBIT_IN32_63 MUX1_1_0 ( .port0({\s_mux1_signals[1][0][31] , 
        \s_mux1_signals[1][0][30] , \s_mux1_signals[1][0][29] , 
        \s_mux1_signals[1][0][28] , \s_mux1_signals[1][0][27] , 
        \s_mux1_signals[1][0][26] , \s_mux1_signals[1][0][25] , 
        \s_mux1_signals[1][0][24] , \s_mux1_signals[1][0][23] , 
        \s_mux1_signals[1][0][22] , \s_mux1_signals[1][0][21] , 
        \s_mux1_signals[1][0][20] , \s_mux1_signals[1][0][19] , 
        \s_mux1_signals[1][0][18] , \s_mux1_signals[1][0][17] , 
        \s_mux1_signals[1][0][16] , \s_mux1_signals[1][0][15] , 
        \s_mux1_signals[1][0][14] , \s_mux1_signals[1][0][13] , 
        \s_mux1_signals[1][0][12] , \s_mux1_signals[1][0][11] , 
        \s_mux1_signals[1][0][10] , \s_mux1_signals[1][0][9] , 
        \s_mux1_signals[1][0][8] , \s_mux1_signals[1][0][7] , 
        \s_mux1_signals[1][0][6] , \s_mux1_signals[1][0][5] , 
        \s_mux1_signals[1][0][4] , \s_mux1_signals[1][0][3] , 
        \s_mux1_signals[1][0][2] , \s_mux1_signals[1][0][1] , 
        \s_mux1_signals[1][0][0] }), .port1({\s_mux1_signals[1][2][31] , 
        \s_mux1_signals[1][2][30] , \s_mux1_signals[1][2][29] , 
        \s_mux1_signals[1][2][28] , \s_mux1_signals[1][2][27] , 
        \s_mux1_signals[1][2][26] , \s_mux1_signals[1][2][25] , 
        \s_mux1_signals[1][2][24] , \s_mux1_signals[1][2][23] , 
        \s_mux1_signals[1][2][22] , \s_mux1_signals[1][2][21] , 
        \s_mux1_signals[1][2][20] , \s_mux1_signals[1][2][19] , 
        \s_mux1_signals[1][2][18] , \s_mux1_signals[1][2][17] , 
        \s_mux1_signals[1][2][16] , \s_mux1_signals[1][2][15] , 
        \s_mux1_signals[1][2][14] , \s_mux1_signals[1][2][13] , 
        \s_mux1_signals[1][2][12] , \s_mux1_signals[1][2][11] , 
        \s_mux1_signals[1][2][10] , \s_mux1_signals[1][2][9] , 
        \s_mux1_signals[1][2][8] , \s_mux1_signals[1][2][7] , 
        \s_mux1_signals[1][2][6] , \s_mux1_signals[1][2][5] , 
        \s_mux1_signals[1][2][4] , \s_mux1_signals[1][2][3] , 
        \s_mux1_signals[1][2][2] , \s_mux1_signals[1][2][1] , 
        \s_mux1_signals[1][2][0] }), .sel(n32), .portY({
        \s_mux1_signals[2][0][31] , \s_mux1_signals[2][0][30] , 
        \s_mux1_signals[2][0][29] , \s_mux1_signals[2][0][28] , 
        \s_mux1_signals[2][0][27] , \s_mux1_signals[2][0][26] , 
        \s_mux1_signals[2][0][25] , \s_mux1_signals[2][0][24] , 
        \s_mux1_signals[2][0][23] , \s_mux1_signals[2][0][22] , 
        \s_mux1_signals[2][0][21] , \s_mux1_signals[2][0][20] , 
        \s_mux1_signals[2][0][19] , \s_mux1_signals[2][0][18] , 
        \s_mux1_signals[2][0][17] , \s_mux1_signals[2][0][16] , 
        \s_mux1_signals[2][0][15] , \s_mux1_signals[2][0][14] , 
        \s_mux1_signals[2][0][13] , \s_mux1_signals[2][0][12] , 
        \s_mux1_signals[2][0][11] , \s_mux1_signals[2][0][10] , 
        \s_mux1_signals[2][0][9] , \s_mux1_signals[2][0][8] , 
        \s_mux1_signals[2][0][7] , \s_mux1_signals[2][0][6] , 
        \s_mux1_signals[2][0][5] , \s_mux1_signals[2][0][4] , 
        \s_mux1_signals[2][0][3] , \s_mux1_signals[2][0][2] , 
        \s_mux1_signals[2][0][1] , \s_mux1_signals[2][0][0] }) );
  Mux_NBit_2x1_NBIT_IN32_62 MUX1_1_4 ( .port0({\s_mux1_signals[1][4][31] , 
        \s_mux1_signals[1][4][30] , \s_mux1_signals[1][4][29] , 
        \s_mux1_signals[1][4][28] , \s_mux1_signals[1][4][27] , 
        \s_mux1_signals[1][4][26] , \s_mux1_signals[1][4][25] , 
        \s_mux1_signals[1][4][24] , \s_mux1_signals[1][4][23] , 
        \s_mux1_signals[1][4][22] , \s_mux1_signals[1][4][21] , 
        \s_mux1_signals[1][4][20] , \s_mux1_signals[1][4][19] , 
        \s_mux1_signals[1][4][18] , \s_mux1_signals[1][4][17] , 
        \s_mux1_signals[1][4][16] , \s_mux1_signals[1][4][15] , 
        \s_mux1_signals[1][4][14] , \s_mux1_signals[1][4][13] , 
        \s_mux1_signals[1][4][12] , \s_mux1_signals[1][4][11] , 
        \s_mux1_signals[1][4][10] , \s_mux1_signals[1][4][9] , 
        \s_mux1_signals[1][4][8] , \s_mux1_signals[1][4][7] , 
        \s_mux1_signals[1][4][6] , \s_mux1_signals[1][4][5] , 
        \s_mux1_signals[1][4][4] , \s_mux1_signals[1][4][3] , 
        \s_mux1_signals[1][4][2] , \s_mux1_signals[1][4][1] , 
        \s_mux1_signals[1][4][0] }), .port1({\s_mux1_signals[1][6][31] , 
        \s_mux1_signals[1][6][30] , \s_mux1_signals[1][6][29] , 
        \s_mux1_signals[1][6][28] , \s_mux1_signals[1][6][27] , 
        \s_mux1_signals[1][6][26] , \s_mux1_signals[1][6][25] , 
        \s_mux1_signals[1][6][24] , \s_mux1_signals[1][6][23] , 
        \s_mux1_signals[1][6][22] , \s_mux1_signals[1][6][21] , 
        \s_mux1_signals[1][6][20] , \s_mux1_signals[1][6][19] , 
        \s_mux1_signals[1][6][18] , \s_mux1_signals[1][6][17] , 
        \s_mux1_signals[1][6][16] , \s_mux1_signals[1][6][15] , 
        \s_mux1_signals[1][6][14] , \s_mux1_signals[1][6][13] , 
        \s_mux1_signals[1][6][12] , \s_mux1_signals[1][6][11] , 
        \s_mux1_signals[1][6][10] , \s_mux1_signals[1][6][9] , 
        \s_mux1_signals[1][6][8] , \s_mux1_signals[1][6][7] , 
        \s_mux1_signals[1][6][6] , \s_mux1_signals[1][6][5] , 
        \s_mux1_signals[1][6][4] , \s_mux1_signals[1][6][3] , 
        \s_mux1_signals[1][6][2] , \s_mux1_signals[1][6][1] , 
        \s_mux1_signals[1][6][0] }), .sel(n32), .portY({
        \s_mux1_signals[2][4][31] , \s_mux1_signals[2][4][30] , 
        \s_mux1_signals[2][4][29] , \s_mux1_signals[2][4][28] , 
        \s_mux1_signals[2][4][27] , \s_mux1_signals[2][4][26] , 
        \s_mux1_signals[2][4][25] , \s_mux1_signals[2][4][24] , 
        \s_mux1_signals[2][4][23] , \s_mux1_signals[2][4][22] , 
        \s_mux1_signals[2][4][21] , \s_mux1_signals[2][4][20] , 
        \s_mux1_signals[2][4][19] , \s_mux1_signals[2][4][18] , 
        \s_mux1_signals[2][4][17] , \s_mux1_signals[2][4][16] , 
        \s_mux1_signals[2][4][15] , \s_mux1_signals[2][4][14] , 
        \s_mux1_signals[2][4][13] , \s_mux1_signals[2][4][12] , 
        \s_mux1_signals[2][4][11] , \s_mux1_signals[2][4][10] , 
        \s_mux1_signals[2][4][9] , \s_mux1_signals[2][4][8] , 
        \s_mux1_signals[2][4][7] , \s_mux1_signals[2][4][6] , 
        \s_mux1_signals[2][4][5] , \s_mux1_signals[2][4][4] , 
        \s_mux1_signals[2][4][3] , \s_mux1_signals[2][4][2] , 
        \s_mux1_signals[2][4][1] , \s_mux1_signals[2][4][0] }) );
  Mux_NBit_2x1_NBIT_IN32_61 MUX1_1_8 ( .port0({\s_mux1_signals[1][8][31] , 
        \s_mux1_signals[1][8][30] , \s_mux1_signals[1][8][29] , 
        \s_mux1_signals[1][8][28] , \s_mux1_signals[1][8][27] , 
        \s_mux1_signals[1][8][26] , \s_mux1_signals[1][8][25] , 
        \s_mux1_signals[1][8][24] , \s_mux1_signals[1][8][23] , 
        \s_mux1_signals[1][8][22] , \s_mux1_signals[1][8][21] , 
        \s_mux1_signals[1][8][20] , \s_mux1_signals[1][8][19] , 
        \s_mux1_signals[1][8][18] , \s_mux1_signals[1][8][17] , 
        \s_mux1_signals[1][8][16] , \s_mux1_signals[1][8][15] , 
        \s_mux1_signals[1][8][14] , \s_mux1_signals[1][8][13] , 
        \s_mux1_signals[1][8][12] , \s_mux1_signals[1][8][11] , 
        \s_mux1_signals[1][8][10] , \s_mux1_signals[1][8][9] , 
        \s_mux1_signals[1][8][8] , \s_mux1_signals[1][8][7] , 
        \s_mux1_signals[1][8][6] , \s_mux1_signals[1][8][5] , 
        \s_mux1_signals[1][8][4] , \s_mux1_signals[1][8][3] , 
        \s_mux1_signals[1][8][2] , \s_mux1_signals[1][8][1] , 
        \s_mux1_signals[1][8][0] }), .port1({\s_mux1_signals[1][10][31] , 
        \s_mux1_signals[1][10][30] , \s_mux1_signals[1][10][29] , 
        \s_mux1_signals[1][10][28] , \s_mux1_signals[1][10][27] , 
        \s_mux1_signals[1][10][26] , \s_mux1_signals[1][10][25] , 
        \s_mux1_signals[1][10][24] , \s_mux1_signals[1][10][23] , 
        \s_mux1_signals[1][10][22] , \s_mux1_signals[1][10][21] , 
        \s_mux1_signals[1][10][20] , \s_mux1_signals[1][10][19] , 
        \s_mux1_signals[1][10][18] , \s_mux1_signals[1][10][17] , 
        \s_mux1_signals[1][10][16] , \s_mux1_signals[1][10][15] , 
        \s_mux1_signals[1][10][14] , \s_mux1_signals[1][10][13] , 
        \s_mux1_signals[1][10][12] , \s_mux1_signals[1][10][11] , 
        \s_mux1_signals[1][10][10] , \s_mux1_signals[1][10][9] , 
        \s_mux1_signals[1][10][8] , \s_mux1_signals[1][10][7] , 
        \s_mux1_signals[1][10][6] , \s_mux1_signals[1][10][5] , 
        \s_mux1_signals[1][10][4] , \s_mux1_signals[1][10][3] , 
        \s_mux1_signals[1][10][2] , \s_mux1_signals[1][10][1] , 
        \s_mux1_signals[1][10][0] }), .sel(n32), .portY({
        \s_mux1_signals[2][8][31] , \s_mux1_signals[2][8][30] , 
        \s_mux1_signals[2][8][29] , \s_mux1_signals[2][8][28] , 
        \s_mux1_signals[2][8][27] , \s_mux1_signals[2][8][26] , 
        \s_mux1_signals[2][8][25] , \s_mux1_signals[2][8][24] , 
        \s_mux1_signals[2][8][23] , \s_mux1_signals[2][8][22] , 
        \s_mux1_signals[2][8][21] , \s_mux1_signals[2][8][20] , 
        \s_mux1_signals[2][8][19] , \s_mux1_signals[2][8][18] , 
        \s_mux1_signals[2][8][17] , \s_mux1_signals[2][8][16] , 
        \s_mux1_signals[2][8][15] , \s_mux1_signals[2][8][14] , 
        \s_mux1_signals[2][8][13] , \s_mux1_signals[2][8][12] , 
        \s_mux1_signals[2][8][11] , \s_mux1_signals[2][8][10] , 
        \s_mux1_signals[2][8][9] , \s_mux1_signals[2][8][8] , 
        \s_mux1_signals[2][8][7] , \s_mux1_signals[2][8][6] , 
        \s_mux1_signals[2][8][5] , \s_mux1_signals[2][8][4] , 
        \s_mux1_signals[2][8][3] , \s_mux1_signals[2][8][2] , 
        \s_mux1_signals[2][8][1] , \s_mux1_signals[2][8][0] }) );
  Mux_NBit_2x1_NBIT_IN32_60 MUX1_1_12 ( .port0({\s_mux1_signals[1][12][31] , 
        \s_mux1_signals[1][12][30] , \s_mux1_signals[1][12][29] , 
        \s_mux1_signals[1][12][28] , \s_mux1_signals[1][12][27] , 
        \s_mux1_signals[1][12][26] , \s_mux1_signals[1][12][25] , 
        \s_mux1_signals[1][12][24] , \s_mux1_signals[1][12][23] , 
        \s_mux1_signals[1][12][22] , \s_mux1_signals[1][12][21] , 
        \s_mux1_signals[1][12][20] , \s_mux1_signals[1][12][19] , 
        \s_mux1_signals[1][12][18] , \s_mux1_signals[1][12][17] , 
        \s_mux1_signals[1][12][16] , \s_mux1_signals[1][12][15] , 
        \s_mux1_signals[1][12][14] , \s_mux1_signals[1][12][13] , 
        \s_mux1_signals[1][12][12] , \s_mux1_signals[1][12][11] , 
        \s_mux1_signals[1][12][10] , \s_mux1_signals[1][12][9] , 
        \s_mux1_signals[1][12][8] , \s_mux1_signals[1][12][7] , 
        \s_mux1_signals[1][12][6] , \s_mux1_signals[1][12][5] , 
        \s_mux1_signals[1][12][4] , \s_mux1_signals[1][12][3] , 
        \s_mux1_signals[1][12][2] , \s_mux1_signals[1][12][1] , 
        \s_mux1_signals[1][12][0] }), .port1({\s_mux1_signals[1][14][31] , 
        \s_mux1_signals[1][14][30] , \s_mux1_signals[1][14][29] , 
        \s_mux1_signals[1][14][28] , \s_mux1_signals[1][14][27] , 
        \s_mux1_signals[1][14][26] , \s_mux1_signals[1][14][25] , 
        \s_mux1_signals[1][14][24] , \s_mux1_signals[1][14][23] , 
        \s_mux1_signals[1][14][22] , \s_mux1_signals[1][14][21] , 
        \s_mux1_signals[1][14][20] , \s_mux1_signals[1][14][19] , 
        \s_mux1_signals[1][14][18] , \s_mux1_signals[1][14][17] , 
        \s_mux1_signals[1][14][16] , \s_mux1_signals[1][14][15] , 
        \s_mux1_signals[1][14][14] , \s_mux1_signals[1][14][13] , 
        \s_mux1_signals[1][14][12] , \s_mux1_signals[1][14][11] , 
        \s_mux1_signals[1][14][10] , \s_mux1_signals[1][14][9] , 
        \s_mux1_signals[1][14][8] , \s_mux1_signals[1][14][7] , 
        \s_mux1_signals[1][14][6] , \s_mux1_signals[1][14][5] , 
        \s_mux1_signals[1][14][4] , \s_mux1_signals[1][14][3] , 
        \s_mux1_signals[1][14][2] , \s_mux1_signals[1][14][1] , 
        \s_mux1_signals[1][14][0] }), .sel(n33), .portY({
        \s_mux1_signals[2][12][31] , \s_mux1_signals[2][12][30] , 
        \s_mux1_signals[2][12][29] , \s_mux1_signals[2][12][28] , 
        \s_mux1_signals[2][12][27] , \s_mux1_signals[2][12][26] , 
        \s_mux1_signals[2][12][25] , \s_mux1_signals[2][12][24] , 
        \s_mux1_signals[2][12][23] , \s_mux1_signals[2][12][22] , 
        \s_mux1_signals[2][12][21] , \s_mux1_signals[2][12][20] , 
        \s_mux1_signals[2][12][19] , \s_mux1_signals[2][12][18] , 
        \s_mux1_signals[2][12][17] , \s_mux1_signals[2][12][16] , 
        \s_mux1_signals[2][12][15] , \s_mux1_signals[2][12][14] , 
        \s_mux1_signals[2][12][13] , \s_mux1_signals[2][12][12] , 
        \s_mux1_signals[2][12][11] , \s_mux1_signals[2][12][10] , 
        \s_mux1_signals[2][12][9] , \s_mux1_signals[2][12][8] , 
        \s_mux1_signals[2][12][7] , \s_mux1_signals[2][12][6] , 
        \s_mux1_signals[2][12][5] , \s_mux1_signals[2][12][4] , 
        \s_mux1_signals[2][12][3] , \s_mux1_signals[2][12][2] , 
        \s_mux1_signals[2][12][1] , \s_mux1_signals[2][12][0] }) );
  Mux_NBit_2x1_NBIT_IN32_59 MUX1_1_16 ( .port0({\s_mux1_signals[1][16][31] , 
        \s_mux1_signals[1][16][30] , \s_mux1_signals[1][16][29] , 
        \s_mux1_signals[1][16][28] , \s_mux1_signals[1][16][27] , 
        \s_mux1_signals[1][16][26] , \s_mux1_signals[1][16][25] , 
        \s_mux1_signals[1][16][24] , \s_mux1_signals[1][16][23] , 
        \s_mux1_signals[1][16][22] , \s_mux1_signals[1][16][21] , 
        \s_mux1_signals[1][16][20] , \s_mux1_signals[1][16][19] , 
        \s_mux1_signals[1][16][18] , \s_mux1_signals[1][16][17] , 
        \s_mux1_signals[1][16][16] , \s_mux1_signals[1][16][15] , 
        \s_mux1_signals[1][16][14] , \s_mux1_signals[1][16][13] , 
        \s_mux1_signals[1][16][12] , \s_mux1_signals[1][16][11] , 
        \s_mux1_signals[1][16][10] , \s_mux1_signals[1][16][9] , 
        \s_mux1_signals[1][16][8] , \s_mux1_signals[1][16][7] , 
        \s_mux1_signals[1][16][6] , \s_mux1_signals[1][16][5] , 
        \s_mux1_signals[1][16][4] , \s_mux1_signals[1][16][3] , 
        \s_mux1_signals[1][16][2] , \s_mux1_signals[1][16][1] , 
        \s_mux1_signals[1][16][0] }), .port1({\s_mux1_signals[1][18][31] , 
        \s_mux1_signals[1][18][30] , \s_mux1_signals[1][18][29] , 
        \s_mux1_signals[1][18][28] , \s_mux1_signals[1][18][27] , 
        \s_mux1_signals[1][18][26] , \s_mux1_signals[1][18][25] , 
        \s_mux1_signals[1][18][24] , \s_mux1_signals[1][18][23] , 
        \s_mux1_signals[1][18][22] , \s_mux1_signals[1][18][21] , 
        \s_mux1_signals[1][18][20] , \s_mux1_signals[1][18][19] , 
        \s_mux1_signals[1][18][18] , \s_mux1_signals[1][18][17] , 
        \s_mux1_signals[1][18][16] , \s_mux1_signals[1][18][15] , 
        \s_mux1_signals[1][18][14] , \s_mux1_signals[1][18][13] , 
        \s_mux1_signals[1][18][12] , \s_mux1_signals[1][18][11] , 
        \s_mux1_signals[1][18][10] , \s_mux1_signals[1][18][9] , 
        \s_mux1_signals[1][18][8] , \s_mux1_signals[1][18][7] , 
        \s_mux1_signals[1][18][6] , \s_mux1_signals[1][18][5] , 
        \s_mux1_signals[1][18][4] , \s_mux1_signals[1][18][3] , 
        \s_mux1_signals[1][18][2] , \s_mux1_signals[1][18][1] , 
        \s_mux1_signals[1][18][0] }), .sel(n33), .portY({
        \s_mux1_signals[2][16][31] , \s_mux1_signals[2][16][30] , 
        \s_mux1_signals[2][16][29] , \s_mux1_signals[2][16][28] , 
        \s_mux1_signals[2][16][27] , \s_mux1_signals[2][16][26] , 
        \s_mux1_signals[2][16][25] , \s_mux1_signals[2][16][24] , 
        \s_mux1_signals[2][16][23] , \s_mux1_signals[2][16][22] , 
        \s_mux1_signals[2][16][21] , \s_mux1_signals[2][16][20] , 
        \s_mux1_signals[2][16][19] , \s_mux1_signals[2][16][18] , 
        \s_mux1_signals[2][16][17] , \s_mux1_signals[2][16][16] , 
        \s_mux1_signals[2][16][15] , \s_mux1_signals[2][16][14] , 
        \s_mux1_signals[2][16][13] , \s_mux1_signals[2][16][12] , 
        \s_mux1_signals[2][16][11] , \s_mux1_signals[2][16][10] , 
        \s_mux1_signals[2][16][9] , \s_mux1_signals[2][16][8] , 
        \s_mux1_signals[2][16][7] , \s_mux1_signals[2][16][6] , 
        \s_mux1_signals[2][16][5] , \s_mux1_signals[2][16][4] , 
        \s_mux1_signals[2][16][3] , \s_mux1_signals[2][16][2] , 
        \s_mux1_signals[2][16][1] , \s_mux1_signals[2][16][0] }) );
  Mux_NBit_2x1_NBIT_IN32_58 MUX1_1_20 ( .port0({\s_mux1_signals[1][20][31] , 
        \s_mux1_signals[1][20][30] , \s_mux1_signals[1][20][29] , 
        \s_mux1_signals[1][20][28] , \s_mux1_signals[1][20][27] , 
        \s_mux1_signals[1][20][26] , \s_mux1_signals[1][20][25] , 
        \s_mux1_signals[1][20][24] , \s_mux1_signals[1][20][23] , 
        \s_mux1_signals[1][20][22] , \s_mux1_signals[1][20][21] , 
        \s_mux1_signals[1][20][20] , \s_mux1_signals[1][20][19] , 
        \s_mux1_signals[1][20][18] , \s_mux1_signals[1][20][17] , 
        \s_mux1_signals[1][20][16] , \s_mux1_signals[1][20][15] , 
        \s_mux1_signals[1][20][14] , \s_mux1_signals[1][20][13] , 
        \s_mux1_signals[1][20][12] , \s_mux1_signals[1][20][11] , 
        \s_mux1_signals[1][20][10] , \s_mux1_signals[1][20][9] , 
        \s_mux1_signals[1][20][8] , \s_mux1_signals[1][20][7] , 
        \s_mux1_signals[1][20][6] , \s_mux1_signals[1][20][5] , 
        \s_mux1_signals[1][20][4] , \s_mux1_signals[1][20][3] , 
        \s_mux1_signals[1][20][2] , \s_mux1_signals[1][20][1] , 
        \s_mux1_signals[1][20][0] }), .port1({\s_mux1_signals[1][22][31] , 
        \s_mux1_signals[1][22][30] , \s_mux1_signals[1][22][29] , 
        \s_mux1_signals[1][22][28] , \s_mux1_signals[1][22][27] , 
        \s_mux1_signals[1][22][26] , \s_mux1_signals[1][22][25] , 
        \s_mux1_signals[1][22][24] , \s_mux1_signals[1][22][23] , 
        \s_mux1_signals[1][22][22] , \s_mux1_signals[1][22][21] , 
        \s_mux1_signals[1][22][20] , \s_mux1_signals[1][22][19] , 
        \s_mux1_signals[1][22][18] , \s_mux1_signals[1][22][17] , 
        \s_mux1_signals[1][22][16] , \s_mux1_signals[1][22][15] , 
        \s_mux1_signals[1][22][14] , \s_mux1_signals[1][22][13] , 
        \s_mux1_signals[1][22][12] , \s_mux1_signals[1][22][11] , 
        \s_mux1_signals[1][22][10] , \s_mux1_signals[1][22][9] , 
        \s_mux1_signals[1][22][8] , \s_mux1_signals[1][22][7] , 
        \s_mux1_signals[1][22][6] , \s_mux1_signals[1][22][5] , 
        \s_mux1_signals[1][22][4] , \s_mux1_signals[1][22][3] , 
        \s_mux1_signals[1][22][2] , \s_mux1_signals[1][22][1] , 
        \s_mux1_signals[1][22][0] }), .sel(n33), .portY({
        \s_mux1_signals[2][20][31] , \s_mux1_signals[2][20][30] , 
        \s_mux1_signals[2][20][29] , \s_mux1_signals[2][20][28] , 
        \s_mux1_signals[2][20][27] , \s_mux1_signals[2][20][26] , 
        \s_mux1_signals[2][20][25] , \s_mux1_signals[2][20][24] , 
        \s_mux1_signals[2][20][23] , \s_mux1_signals[2][20][22] , 
        \s_mux1_signals[2][20][21] , \s_mux1_signals[2][20][20] , 
        \s_mux1_signals[2][20][19] , \s_mux1_signals[2][20][18] , 
        \s_mux1_signals[2][20][17] , \s_mux1_signals[2][20][16] , 
        \s_mux1_signals[2][20][15] , \s_mux1_signals[2][20][14] , 
        \s_mux1_signals[2][20][13] , \s_mux1_signals[2][20][12] , 
        \s_mux1_signals[2][20][11] , \s_mux1_signals[2][20][10] , 
        \s_mux1_signals[2][20][9] , \s_mux1_signals[2][20][8] , 
        \s_mux1_signals[2][20][7] , \s_mux1_signals[2][20][6] , 
        \s_mux1_signals[2][20][5] , \s_mux1_signals[2][20][4] , 
        \s_mux1_signals[2][20][3] , \s_mux1_signals[2][20][2] , 
        \s_mux1_signals[2][20][1] , \s_mux1_signals[2][20][0] }) );
  Mux_NBit_2x1_NBIT_IN32_57 MUX1_1_24 ( .port0({\s_mux1_signals[1][24][31] , 
        \s_mux1_signals[1][24][30] , \s_mux1_signals[1][24][29] , 
        \s_mux1_signals[1][24][28] , \s_mux1_signals[1][24][27] , 
        \s_mux1_signals[1][24][26] , \s_mux1_signals[1][24][25] , 
        \s_mux1_signals[1][24][24] , \s_mux1_signals[1][24][23] , 
        \s_mux1_signals[1][24][22] , \s_mux1_signals[1][24][21] , 
        \s_mux1_signals[1][24][20] , \s_mux1_signals[1][24][19] , 
        \s_mux1_signals[1][24][18] , \s_mux1_signals[1][24][17] , 
        \s_mux1_signals[1][24][16] , \s_mux1_signals[1][24][15] , 
        \s_mux1_signals[1][24][14] , \s_mux1_signals[1][24][13] , 
        \s_mux1_signals[1][24][12] , \s_mux1_signals[1][24][11] , 
        \s_mux1_signals[1][24][10] , \s_mux1_signals[1][24][9] , 
        \s_mux1_signals[1][24][8] , \s_mux1_signals[1][24][7] , 
        \s_mux1_signals[1][24][6] , \s_mux1_signals[1][24][5] , 
        \s_mux1_signals[1][24][4] , \s_mux1_signals[1][24][3] , 
        \s_mux1_signals[1][24][2] , \s_mux1_signals[1][24][1] , 
        \s_mux1_signals[1][24][0] }), .port1({\s_mux1_signals[1][26][31] , 
        \s_mux1_signals[1][26][30] , \s_mux1_signals[1][26][29] , 
        \s_mux1_signals[1][26][28] , \s_mux1_signals[1][26][27] , 
        \s_mux1_signals[1][26][26] , \s_mux1_signals[1][26][25] , 
        \s_mux1_signals[1][26][24] , \s_mux1_signals[1][26][23] , 
        \s_mux1_signals[1][26][22] , \s_mux1_signals[1][26][21] , 
        \s_mux1_signals[1][26][20] , \s_mux1_signals[1][26][19] , 
        \s_mux1_signals[1][26][18] , \s_mux1_signals[1][26][17] , 
        \s_mux1_signals[1][26][16] , \s_mux1_signals[1][26][15] , 
        \s_mux1_signals[1][26][14] , \s_mux1_signals[1][26][13] , 
        \s_mux1_signals[1][26][12] , \s_mux1_signals[1][26][11] , 
        \s_mux1_signals[1][26][10] , \s_mux1_signals[1][26][9] , 
        \s_mux1_signals[1][26][8] , \s_mux1_signals[1][26][7] , 
        \s_mux1_signals[1][26][6] , \s_mux1_signals[1][26][5] , 
        \s_mux1_signals[1][26][4] , \s_mux1_signals[1][26][3] , 
        \s_mux1_signals[1][26][2] , \s_mux1_signals[1][26][1] , 
        \s_mux1_signals[1][26][0] }), .sel(n34), .portY({
        \s_mux1_signals[2][24][31] , \s_mux1_signals[2][24][30] , 
        \s_mux1_signals[2][24][29] , \s_mux1_signals[2][24][28] , 
        \s_mux1_signals[2][24][27] , \s_mux1_signals[2][24][26] , 
        \s_mux1_signals[2][24][25] , \s_mux1_signals[2][24][24] , 
        \s_mux1_signals[2][24][23] , \s_mux1_signals[2][24][22] , 
        \s_mux1_signals[2][24][21] , \s_mux1_signals[2][24][20] , 
        \s_mux1_signals[2][24][19] , \s_mux1_signals[2][24][18] , 
        \s_mux1_signals[2][24][17] , \s_mux1_signals[2][24][16] , 
        \s_mux1_signals[2][24][15] , \s_mux1_signals[2][24][14] , 
        \s_mux1_signals[2][24][13] , \s_mux1_signals[2][24][12] , 
        \s_mux1_signals[2][24][11] , \s_mux1_signals[2][24][10] , 
        \s_mux1_signals[2][24][9] , \s_mux1_signals[2][24][8] , 
        \s_mux1_signals[2][24][7] , \s_mux1_signals[2][24][6] , 
        \s_mux1_signals[2][24][5] , \s_mux1_signals[2][24][4] , 
        \s_mux1_signals[2][24][3] , \s_mux1_signals[2][24][2] , 
        \s_mux1_signals[2][24][1] , \s_mux1_signals[2][24][0] }) );
  Mux_NBit_2x1_NBIT_IN32_56 MUX1_1_28 ( .port0({\s_mux1_signals[1][28][31] , 
        \s_mux1_signals[1][28][30] , \s_mux1_signals[1][28][29] , 
        \s_mux1_signals[1][28][28] , \s_mux1_signals[1][28][27] , 
        \s_mux1_signals[1][28][26] , \s_mux1_signals[1][28][25] , 
        \s_mux1_signals[1][28][24] , \s_mux1_signals[1][28][23] , 
        \s_mux1_signals[1][28][22] , \s_mux1_signals[1][28][21] , 
        \s_mux1_signals[1][28][20] , \s_mux1_signals[1][28][19] , 
        \s_mux1_signals[1][28][18] , \s_mux1_signals[1][28][17] , 
        \s_mux1_signals[1][28][16] , \s_mux1_signals[1][28][15] , 
        \s_mux1_signals[1][28][14] , \s_mux1_signals[1][28][13] , 
        \s_mux1_signals[1][28][12] , \s_mux1_signals[1][28][11] , 
        \s_mux1_signals[1][28][10] , \s_mux1_signals[1][28][9] , 
        \s_mux1_signals[1][28][8] , \s_mux1_signals[1][28][7] , 
        \s_mux1_signals[1][28][6] , \s_mux1_signals[1][28][5] , 
        \s_mux1_signals[1][28][4] , \s_mux1_signals[1][28][3] , 
        \s_mux1_signals[1][28][2] , \s_mux1_signals[1][28][1] , 
        \s_mux1_signals[1][28][0] }), .port1({\s_mux1_signals[1][30][31] , 
        \s_mux1_signals[1][30][30] , \s_mux1_signals[1][30][29] , 
        \s_mux1_signals[1][30][28] , \s_mux1_signals[1][30][27] , 
        \s_mux1_signals[1][30][26] , \s_mux1_signals[1][30][25] , 
        \s_mux1_signals[1][30][24] , \s_mux1_signals[1][30][23] , 
        \s_mux1_signals[1][30][22] , \s_mux1_signals[1][30][21] , 
        \s_mux1_signals[1][30][20] , \s_mux1_signals[1][30][19] , 
        \s_mux1_signals[1][30][18] , \s_mux1_signals[1][30][17] , 
        \s_mux1_signals[1][30][16] , \s_mux1_signals[1][30][15] , 
        \s_mux1_signals[1][30][14] , \s_mux1_signals[1][30][13] , 
        \s_mux1_signals[1][30][12] , \s_mux1_signals[1][30][11] , 
        \s_mux1_signals[1][30][10] , \s_mux1_signals[1][30][9] , 
        \s_mux1_signals[1][30][8] , \s_mux1_signals[1][30][7] , 
        \s_mux1_signals[1][30][6] , \s_mux1_signals[1][30][5] , 
        \s_mux1_signals[1][30][4] , \s_mux1_signals[1][30][3] , 
        \s_mux1_signals[1][30][2] , \s_mux1_signals[1][30][1] , 
        \s_mux1_signals[1][30][0] }), .sel(n34), .portY({
        \s_mux1_signals[2][28][31] , \s_mux1_signals[2][28][30] , 
        \s_mux1_signals[2][28][29] , \s_mux1_signals[2][28][28] , 
        \s_mux1_signals[2][28][27] , \s_mux1_signals[2][28][26] , 
        \s_mux1_signals[2][28][25] , \s_mux1_signals[2][28][24] , 
        \s_mux1_signals[2][28][23] , \s_mux1_signals[2][28][22] , 
        \s_mux1_signals[2][28][21] , \s_mux1_signals[2][28][20] , 
        \s_mux1_signals[2][28][19] , \s_mux1_signals[2][28][18] , 
        \s_mux1_signals[2][28][17] , \s_mux1_signals[2][28][16] , 
        \s_mux1_signals[2][28][15] , \s_mux1_signals[2][28][14] , 
        \s_mux1_signals[2][28][13] , \s_mux1_signals[2][28][12] , 
        \s_mux1_signals[2][28][11] , \s_mux1_signals[2][28][10] , 
        \s_mux1_signals[2][28][9] , \s_mux1_signals[2][28][8] , 
        \s_mux1_signals[2][28][7] , \s_mux1_signals[2][28][6] , 
        \s_mux1_signals[2][28][5] , \s_mux1_signals[2][28][4] , 
        \s_mux1_signals[2][28][3] , \s_mux1_signals[2][28][2] , 
        \s_mux1_signals[2][28][1] , \s_mux1_signals[2][28][0] }) );
  Mux_NBit_2x1_NBIT_IN32_55 MUX1_2_0 ( .port0({\s_mux1_signals[2][0][31] , 
        \s_mux1_signals[2][0][30] , \s_mux1_signals[2][0][29] , 
        \s_mux1_signals[2][0][28] , \s_mux1_signals[2][0][27] , 
        \s_mux1_signals[2][0][26] , \s_mux1_signals[2][0][25] , 
        \s_mux1_signals[2][0][24] , \s_mux1_signals[2][0][23] , 
        \s_mux1_signals[2][0][22] , \s_mux1_signals[2][0][21] , 
        \s_mux1_signals[2][0][20] , \s_mux1_signals[2][0][19] , 
        \s_mux1_signals[2][0][18] , \s_mux1_signals[2][0][17] , 
        \s_mux1_signals[2][0][16] , \s_mux1_signals[2][0][15] , 
        \s_mux1_signals[2][0][14] , \s_mux1_signals[2][0][13] , 
        \s_mux1_signals[2][0][12] , \s_mux1_signals[2][0][11] , 
        \s_mux1_signals[2][0][10] , \s_mux1_signals[2][0][9] , 
        \s_mux1_signals[2][0][8] , \s_mux1_signals[2][0][7] , 
        \s_mux1_signals[2][0][6] , \s_mux1_signals[2][0][5] , 
        \s_mux1_signals[2][0][4] , \s_mux1_signals[2][0][3] , 
        \s_mux1_signals[2][0][2] , \s_mux1_signals[2][0][1] , 
        \s_mux1_signals[2][0][0] }), .port1({\s_mux1_signals[2][4][31] , 
        \s_mux1_signals[2][4][30] , \s_mux1_signals[2][4][29] , 
        \s_mux1_signals[2][4][28] , \s_mux1_signals[2][4][27] , 
        \s_mux1_signals[2][4][26] , \s_mux1_signals[2][4][25] , 
        \s_mux1_signals[2][4][24] , \s_mux1_signals[2][4][23] , 
        \s_mux1_signals[2][4][22] , \s_mux1_signals[2][4][21] , 
        \s_mux1_signals[2][4][20] , \s_mux1_signals[2][4][19] , 
        \s_mux1_signals[2][4][18] , \s_mux1_signals[2][4][17] , 
        \s_mux1_signals[2][4][16] , \s_mux1_signals[2][4][15] , 
        \s_mux1_signals[2][4][14] , \s_mux1_signals[2][4][13] , 
        \s_mux1_signals[2][4][12] , \s_mux1_signals[2][4][11] , 
        \s_mux1_signals[2][4][10] , \s_mux1_signals[2][4][9] , 
        \s_mux1_signals[2][4][8] , \s_mux1_signals[2][4][7] , 
        \s_mux1_signals[2][4][6] , \s_mux1_signals[2][4][5] , 
        \s_mux1_signals[2][4][4] , \s_mux1_signals[2][4][3] , 
        \s_mux1_signals[2][4][2] , \s_mux1_signals[2][4][1] , 
        \s_mux1_signals[2][4][0] }), .sel(n35), .portY({
        \s_mux1_signals[3][0][31] , \s_mux1_signals[3][0][30] , 
        \s_mux1_signals[3][0][29] , \s_mux1_signals[3][0][28] , 
        \s_mux1_signals[3][0][27] , \s_mux1_signals[3][0][26] , 
        \s_mux1_signals[3][0][25] , \s_mux1_signals[3][0][24] , 
        \s_mux1_signals[3][0][23] , \s_mux1_signals[3][0][22] , 
        \s_mux1_signals[3][0][21] , \s_mux1_signals[3][0][20] , 
        \s_mux1_signals[3][0][19] , \s_mux1_signals[3][0][18] , 
        \s_mux1_signals[3][0][17] , \s_mux1_signals[3][0][16] , 
        \s_mux1_signals[3][0][15] , \s_mux1_signals[3][0][14] , 
        \s_mux1_signals[3][0][13] , \s_mux1_signals[3][0][12] , 
        \s_mux1_signals[3][0][11] , \s_mux1_signals[3][0][10] , 
        \s_mux1_signals[3][0][9] , \s_mux1_signals[3][0][8] , 
        \s_mux1_signals[3][0][7] , \s_mux1_signals[3][0][6] , 
        \s_mux1_signals[3][0][5] , \s_mux1_signals[3][0][4] , 
        \s_mux1_signals[3][0][3] , \s_mux1_signals[3][0][2] , 
        \s_mux1_signals[3][0][1] , \s_mux1_signals[3][0][0] }) );
  Mux_NBit_2x1_NBIT_IN32_54 MUX1_2_8 ( .port0({\s_mux1_signals[2][8][31] , 
        \s_mux1_signals[2][8][30] , \s_mux1_signals[2][8][29] , 
        \s_mux1_signals[2][8][28] , \s_mux1_signals[2][8][27] , 
        \s_mux1_signals[2][8][26] , \s_mux1_signals[2][8][25] , 
        \s_mux1_signals[2][8][24] , \s_mux1_signals[2][8][23] , 
        \s_mux1_signals[2][8][22] , \s_mux1_signals[2][8][21] , 
        \s_mux1_signals[2][8][20] , \s_mux1_signals[2][8][19] , 
        \s_mux1_signals[2][8][18] , \s_mux1_signals[2][8][17] , 
        \s_mux1_signals[2][8][16] , \s_mux1_signals[2][8][15] , 
        \s_mux1_signals[2][8][14] , \s_mux1_signals[2][8][13] , 
        \s_mux1_signals[2][8][12] , \s_mux1_signals[2][8][11] , 
        \s_mux1_signals[2][8][10] , \s_mux1_signals[2][8][9] , 
        \s_mux1_signals[2][8][8] , \s_mux1_signals[2][8][7] , 
        \s_mux1_signals[2][8][6] , \s_mux1_signals[2][8][5] , 
        \s_mux1_signals[2][8][4] , \s_mux1_signals[2][8][3] , 
        \s_mux1_signals[2][8][2] , \s_mux1_signals[2][8][1] , 
        \s_mux1_signals[2][8][0] }), .port1({\s_mux1_signals[2][12][31] , 
        \s_mux1_signals[2][12][30] , \s_mux1_signals[2][12][29] , 
        \s_mux1_signals[2][12][28] , \s_mux1_signals[2][12][27] , 
        \s_mux1_signals[2][12][26] , \s_mux1_signals[2][12][25] , 
        \s_mux1_signals[2][12][24] , \s_mux1_signals[2][12][23] , 
        \s_mux1_signals[2][12][22] , \s_mux1_signals[2][12][21] , 
        \s_mux1_signals[2][12][20] , \s_mux1_signals[2][12][19] , 
        \s_mux1_signals[2][12][18] , \s_mux1_signals[2][12][17] , 
        \s_mux1_signals[2][12][16] , \s_mux1_signals[2][12][15] , 
        \s_mux1_signals[2][12][14] , \s_mux1_signals[2][12][13] , 
        \s_mux1_signals[2][12][12] , \s_mux1_signals[2][12][11] , 
        \s_mux1_signals[2][12][10] , \s_mux1_signals[2][12][9] , 
        \s_mux1_signals[2][12][8] , \s_mux1_signals[2][12][7] , 
        \s_mux1_signals[2][12][6] , \s_mux1_signals[2][12][5] , 
        \s_mux1_signals[2][12][4] , \s_mux1_signals[2][12][3] , 
        \s_mux1_signals[2][12][2] , \s_mux1_signals[2][12][1] , 
        \s_mux1_signals[2][12][0] }), .sel(n35), .portY({
        \s_mux1_signals[3][8][31] , \s_mux1_signals[3][8][30] , 
        \s_mux1_signals[3][8][29] , \s_mux1_signals[3][8][28] , 
        \s_mux1_signals[3][8][27] , \s_mux1_signals[3][8][26] , 
        \s_mux1_signals[3][8][25] , \s_mux1_signals[3][8][24] , 
        \s_mux1_signals[3][8][23] , \s_mux1_signals[3][8][22] , 
        \s_mux1_signals[3][8][21] , \s_mux1_signals[3][8][20] , 
        \s_mux1_signals[3][8][19] , \s_mux1_signals[3][8][18] , 
        \s_mux1_signals[3][8][17] , \s_mux1_signals[3][8][16] , 
        \s_mux1_signals[3][8][15] , \s_mux1_signals[3][8][14] , 
        \s_mux1_signals[3][8][13] , \s_mux1_signals[3][8][12] , 
        \s_mux1_signals[3][8][11] , \s_mux1_signals[3][8][10] , 
        \s_mux1_signals[3][8][9] , \s_mux1_signals[3][8][8] , 
        \s_mux1_signals[3][8][7] , \s_mux1_signals[3][8][6] , 
        \s_mux1_signals[3][8][5] , \s_mux1_signals[3][8][4] , 
        \s_mux1_signals[3][8][3] , \s_mux1_signals[3][8][2] , 
        \s_mux1_signals[3][8][1] , \s_mux1_signals[3][8][0] }) );
  Mux_NBit_2x1_NBIT_IN32_53 MUX1_2_16 ( .port0({\s_mux1_signals[2][16][31] , 
        \s_mux1_signals[2][16][30] , \s_mux1_signals[2][16][29] , 
        \s_mux1_signals[2][16][28] , \s_mux1_signals[2][16][27] , 
        \s_mux1_signals[2][16][26] , \s_mux1_signals[2][16][25] , 
        \s_mux1_signals[2][16][24] , \s_mux1_signals[2][16][23] , 
        \s_mux1_signals[2][16][22] , \s_mux1_signals[2][16][21] , 
        \s_mux1_signals[2][16][20] , \s_mux1_signals[2][16][19] , 
        \s_mux1_signals[2][16][18] , \s_mux1_signals[2][16][17] , 
        \s_mux1_signals[2][16][16] , \s_mux1_signals[2][16][15] , 
        \s_mux1_signals[2][16][14] , \s_mux1_signals[2][16][13] , 
        \s_mux1_signals[2][16][12] , \s_mux1_signals[2][16][11] , 
        \s_mux1_signals[2][16][10] , \s_mux1_signals[2][16][9] , 
        \s_mux1_signals[2][16][8] , \s_mux1_signals[2][16][7] , 
        \s_mux1_signals[2][16][6] , \s_mux1_signals[2][16][5] , 
        \s_mux1_signals[2][16][4] , \s_mux1_signals[2][16][3] , 
        \s_mux1_signals[2][16][2] , \s_mux1_signals[2][16][1] , 
        \s_mux1_signals[2][16][0] }), .port1({\s_mux1_signals[2][20][31] , 
        \s_mux1_signals[2][20][30] , \s_mux1_signals[2][20][29] , 
        \s_mux1_signals[2][20][28] , \s_mux1_signals[2][20][27] , 
        \s_mux1_signals[2][20][26] , \s_mux1_signals[2][20][25] , 
        \s_mux1_signals[2][20][24] , \s_mux1_signals[2][20][23] , 
        \s_mux1_signals[2][20][22] , \s_mux1_signals[2][20][21] , 
        \s_mux1_signals[2][20][20] , \s_mux1_signals[2][20][19] , 
        \s_mux1_signals[2][20][18] , \s_mux1_signals[2][20][17] , 
        \s_mux1_signals[2][20][16] , \s_mux1_signals[2][20][15] , 
        \s_mux1_signals[2][20][14] , \s_mux1_signals[2][20][13] , 
        \s_mux1_signals[2][20][12] , \s_mux1_signals[2][20][11] , 
        \s_mux1_signals[2][20][10] , \s_mux1_signals[2][20][9] , 
        \s_mux1_signals[2][20][8] , \s_mux1_signals[2][20][7] , 
        \s_mux1_signals[2][20][6] , \s_mux1_signals[2][20][5] , 
        \s_mux1_signals[2][20][4] , \s_mux1_signals[2][20][3] , 
        \s_mux1_signals[2][20][2] , \s_mux1_signals[2][20][1] , 
        \s_mux1_signals[2][20][0] }), .sel(n35), .portY({
        \s_mux1_signals[3][16][31] , \s_mux1_signals[3][16][30] , 
        \s_mux1_signals[3][16][29] , \s_mux1_signals[3][16][28] , 
        \s_mux1_signals[3][16][27] , \s_mux1_signals[3][16][26] , 
        \s_mux1_signals[3][16][25] , \s_mux1_signals[3][16][24] , 
        \s_mux1_signals[3][16][23] , \s_mux1_signals[3][16][22] , 
        \s_mux1_signals[3][16][21] , \s_mux1_signals[3][16][20] , 
        \s_mux1_signals[3][16][19] , \s_mux1_signals[3][16][18] , 
        \s_mux1_signals[3][16][17] , \s_mux1_signals[3][16][16] , 
        \s_mux1_signals[3][16][15] , \s_mux1_signals[3][16][14] , 
        \s_mux1_signals[3][16][13] , \s_mux1_signals[3][16][12] , 
        \s_mux1_signals[3][16][11] , \s_mux1_signals[3][16][10] , 
        \s_mux1_signals[3][16][9] , \s_mux1_signals[3][16][8] , 
        \s_mux1_signals[3][16][7] , \s_mux1_signals[3][16][6] , 
        \s_mux1_signals[3][16][5] , \s_mux1_signals[3][16][4] , 
        \s_mux1_signals[3][16][3] , \s_mux1_signals[3][16][2] , 
        \s_mux1_signals[3][16][1] , \s_mux1_signals[3][16][0] }) );
  Mux_NBit_2x1_NBIT_IN32_52 MUX1_2_24 ( .port0({\s_mux1_signals[2][24][31] , 
        \s_mux1_signals[2][24][30] , \s_mux1_signals[2][24][29] , 
        \s_mux1_signals[2][24][28] , \s_mux1_signals[2][24][27] , 
        \s_mux1_signals[2][24][26] , \s_mux1_signals[2][24][25] , 
        \s_mux1_signals[2][24][24] , \s_mux1_signals[2][24][23] , 
        \s_mux1_signals[2][24][22] , \s_mux1_signals[2][24][21] , 
        \s_mux1_signals[2][24][20] , \s_mux1_signals[2][24][19] , 
        \s_mux1_signals[2][24][18] , \s_mux1_signals[2][24][17] , 
        \s_mux1_signals[2][24][16] , \s_mux1_signals[2][24][15] , 
        \s_mux1_signals[2][24][14] , \s_mux1_signals[2][24][13] , 
        \s_mux1_signals[2][24][12] , \s_mux1_signals[2][24][11] , 
        \s_mux1_signals[2][24][10] , \s_mux1_signals[2][24][9] , 
        \s_mux1_signals[2][24][8] , \s_mux1_signals[2][24][7] , 
        \s_mux1_signals[2][24][6] , \s_mux1_signals[2][24][5] , 
        \s_mux1_signals[2][24][4] , \s_mux1_signals[2][24][3] , 
        \s_mux1_signals[2][24][2] , \s_mux1_signals[2][24][1] , 
        \s_mux1_signals[2][24][0] }), .port1({\s_mux1_signals[2][28][31] , 
        \s_mux1_signals[2][28][30] , \s_mux1_signals[2][28][29] , 
        \s_mux1_signals[2][28][28] , \s_mux1_signals[2][28][27] , 
        \s_mux1_signals[2][28][26] , \s_mux1_signals[2][28][25] , 
        \s_mux1_signals[2][28][24] , \s_mux1_signals[2][28][23] , 
        \s_mux1_signals[2][28][22] , \s_mux1_signals[2][28][21] , 
        \s_mux1_signals[2][28][20] , \s_mux1_signals[2][28][19] , 
        \s_mux1_signals[2][28][18] , \s_mux1_signals[2][28][17] , 
        \s_mux1_signals[2][28][16] , \s_mux1_signals[2][28][15] , 
        \s_mux1_signals[2][28][14] , \s_mux1_signals[2][28][13] , 
        \s_mux1_signals[2][28][12] , \s_mux1_signals[2][28][11] , 
        \s_mux1_signals[2][28][10] , \s_mux1_signals[2][28][9] , 
        \s_mux1_signals[2][28][8] , \s_mux1_signals[2][28][7] , 
        \s_mux1_signals[2][28][6] , \s_mux1_signals[2][28][5] , 
        \s_mux1_signals[2][28][4] , \s_mux1_signals[2][28][3] , 
        \s_mux1_signals[2][28][2] , \s_mux1_signals[2][28][1] , 
        \s_mux1_signals[2][28][0] }), .sel(n35), .portY({
        \s_mux1_signals[3][24][31] , \s_mux1_signals[3][24][30] , 
        \s_mux1_signals[3][24][29] , \s_mux1_signals[3][24][28] , 
        \s_mux1_signals[3][24][27] , \s_mux1_signals[3][24][26] , 
        \s_mux1_signals[3][24][25] , \s_mux1_signals[3][24][24] , 
        \s_mux1_signals[3][24][23] , \s_mux1_signals[3][24][22] , 
        \s_mux1_signals[3][24][21] , \s_mux1_signals[3][24][20] , 
        \s_mux1_signals[3][24][19] , \s_mux1_signals[3][24][18] , 
        \s_mux1_signals[3][24][17] , \s_mux1_signals[3][24][16] , 
        \s_mux1_signals[3][24][15] , \s_mux1_signals[3][24][14] , 
        \s_mux1_signals[3][24][13] , \s_mux1_signals[3][24][12] , 
        \s_mux1_signals[3][24][11] , \s_mux1_signals[3][24][10] , 
        \s_mux1_signals[3][24][9] , \s_mux1_signals[3][24][8] , 
        \s_mux1_signals[3][24][7] , \s_mux1_signals[3][24][6] , 
        \s_mux1_signals[3][24][5] , \s_mux1_signals[3][24][4] , 
        \s_mux1_signals[3][24][3] , \s_mux1_signals[3][24][2] , 
        \s_mux1_signals[3][24][1] , \s_mux1_signals[3][24][0] }) );
  Mux_NBit_2x1_NBIT_IN32_51 MUX1_3_0 ( .port0({\s_mux1_signals[3][0][31] , 
        \s_mux1_signals[3][0][30] , \s_mux1_signals[3][0][29] , 
        \s_mux1_signals[3][0][28] , \s_mux1_signals[3][0][27] , 
        \s_mux1_signals[3][0][26] , \s_mux1_signals[3][0][25] , 
        \s_mux1_signals[3][0][24] , \s_mux1_signals[3][0][23] , 
        \s_mux1_signals[3][0][22] , \s_mux1_signals[3][0][21] , 
        \s_mux1_signals[3][0][20] , \s_mux1_signals[3][0][19] , 
        \s_mux1_signals[3][0][18] , \s_mux1_signals[3][0][17] , 
        \s_mux1_signals[3][0][16] , \s_mux1_signals[3][0][15] , 
        \s_mux1_signals[3][0][14] , \s_mux1_signals[3][0][13] , 
        \s_mux1_signals[3][0][12] , \s_mux1_signals[3][0][11] , 
        \s_mux1_signals[3][0][10] , \s_mux1_signals[3][0][9] , 
        \s_mux1_signals[3][0][8] , \s_mux1_signals[3][0][7] , 
        \s_mux1_signals[3][0][6] , \s_mux1_signals[3][0][5] , 
        \s_mux1_signals[3][0][4] , \s_mux1_signals[3][0][3] , 
        \s_mux1_signals[3][0][2] , \s_mux1_signals[3][0][1] , 
        \s_mux1_signals[3][0][0] }), .port1({\s_mux1_signals[3][8][31] , 
        \s_mux1_signals[3][8][30] , \s_mux1_signals[3][8][29] , 
        \s_mux1_signals[3][8][28] , \s_mux1_signals[3][8][27] , 
        \s_mux1_signals[3][8][26] , \s_mux1_signals[3][8][25] , 
        \s_mux1_signals[3][8][24] , \s_mux1_signals[3][8][23] , 
        \s_mux1_signals[3][8][22] , \s_mux1_signals[3][8][21] , 
        \s_mux1_signals[3][8][20] , \s_mux1_signals[3][8][19] , 
        \s_mux1_signals[3][8][18] , \s_mux1_signals[3][8][17] , 
        \s_mux1_signals[3][8][16] , \s_mux1_signals[3][8][15] , 
        \s_mux1_signals[3][8][14] , \s_mux1_signals[3][8][13] , 
        \s_mux1_signals[3][8][12] , \s_mux1_signals[3][8][11] , 
        \s_mux1_signals[3][8][10] , \s_mux1_signals[3][8][9] , 
        \s_mux1_signals[3][8][8] , \s_mux1_signals[3][8][7] , 
        \s_mux1_signals[3][8][6] , \s_mux1_signals[3][8][5] , 
        \s_mux1_signals[3][8][4] , \s_mux1_signals[3][8][3] , 
        \s_mux1_signals[3][8][2] , \s_mux1_signals[3][8][1] , 
        \s_mux1_signals[3][8][0] }), .sel(s_addrRd1_Fei_Tmux[3]), .portY({
        \s_mux1_signals[4][0][31] , \s_mux1_signals[4][0][30] , 
        \s_mux1_signals[4][0][29] , \s_mux1_signals[4][0][28] , 
        \s_mux1_signals[4][0][27] , \s_mux1_signals[4][0][26] , 
        \s_mux1_signals[4][0][25] , \s_mux1_signals[4][0][24] , 
        \s_mux1_signals[4][0][23] , \s_mux1_signals[4][0][22] , 
        \s_mux1_signals[4][0][21] , \s_mux1_signals[4][0][20] , 
        \s_mux1_signals[4][0][19] , \s_mux1_signals[4][0][18] , 
        \s_mux1_signals[4][0][17] , \s_mux1_signals[4][0][16] , 
        \s_mux1_signals[4][0][15] , \s_mux1_signals[4][0][14] , 
        \s_mux1_signals[4][0][13] , \s_mux1_signals[4][0][12] , 
        \s_mux1_signals[4][0][11] , \s_mux1_signals[4][0][10] , 
        \s_mux1_signals[4][0][9] , \s_mux1_signals[4][0][8] , 
        \s_mux1_signals[4][0][7] , \s_mux1_signals[4][0][6] , 
        \s_mux1_signals[4][0][5] , \s_mux1_signals[4][0][4] , 
        \s_mux1_signals[4][0][3] , \s_mux1_signals[4][0][2] , 
        \s_mux1_signals[4][0][1] , \s_mux1_signals[4][0][0] }) );
  Mux_NBit_2x1_NBIT_IN32_50 MUX1_3_16 ( .port0({\s_mux1_signals[3][16][31] , 
        \s_mux1_signals[3][16][30] , \s_mux1_signals[3][16][29] , 
        \s_mux1_signals[3][16][28] , \s_mux1_signals[3][16][27] , 
        \s_mux1_signals[3][16][26] , \s_mux1_signals[3][16][25] , 
        \s_mux1_signals[3][16][24] , \s_mux1_signals[3][16][23] , 
        \s_mux1_signals[3][16][22] , \s_mux1_signals[3][16][21] , 
        \s_mux1_signals[3][16][20] , \s_mux1_signals[3][16][19] , 
        \s_mux1_signals[3][16][18] , \s_mux1_signals[3][16][17] , 
        \s_mux1_signals[3][16][16] , \s_mux1_signals[3][16][15] , 
        \s_mux1_signals[3][16][14] , \s_mux1_signals[3][16][13] , 
        \s_mux1_signals[3][16][12] , \s_mux1_signals[3][16][11] , 
        \s_mux1_signals[3][16][10] , \s_mux1_signals[3][16][9] , 
        \s_mux1_signals[3][16][8] , \s_mux1_signals[3][16][7] , 
        \s_mux1_signals[3][16][6] , \s_mux1_signals[3][16][5] , 
        \s_mux1_signals[3][16][4] , \s_mux1_signals[3][16][3] , 
        \s_mux1_signals[3][16][2] , \s_mux1_signals[3][16][1] , 
        \s_mux1_signals[3][16][0] }), .port1({\s_mux1_signals[3][24][31] , 
        \s_mux1_signals[3][24][30] , \s_mux1_signals[3][24][29] , 
        \s_mux1_signals[3][24][28] , \s_mux1_signals[3][24][27] , 
        \s_mux1_signals[3][24][26] , \s_mux1_signals[3][24][25] , 
        \s_mux1_signals[3][24][24] , \s_mux1_signals[3][24][23] , 
        \s_mux1_signals[3][24][22] , \s_mux1_signals[3][24][21] , 
        \s_mux1_signals[3][24][20] , \s_mux1_signals[3][24][19] , 
        \s_mux1_signals[3][24][18] , \s_mux1_signals[3][24][17] , 
        \s_mux1_signals[3][24][16] , \s_mux1_signals[3][24][15] , 
        \s_mux1_signals[3][24][14] , \s_mux1_signals[3][24][13] , 
        \s_mux1_signals[3][24][12] , \s_mux1_signals[3][24][11] , 
        \s_mux1_signals[3][24][10] , \s_mux1_signals[3][24][9] , 
        \s_mux1_signals[3][24][8] , \s_mux1_signals[3][24][7] , 
        \s_mux1_signals[3][24][6] , \s_mux1_signals[3][24][5] , 
        \s_mux1_signals[3][24][4] , \s_mux1_signals[3][24][3] , 
        \s_mux1_signals[3][24][2] , \s_mux1_signals[3][24][1] , 
        \s_mux1_signals[3][24][0] }), .sel(s_addrRd1_Fei_Tmux[3]), .portY({
        \s_mux1_signals[4][16][31] , \s_mux1_signals[4][16][30] , 
        \s_mux1_signals[4][16][29] , \s_mux1_signals[4][16][28] , 
        \s_mux1_signals[4][16][27] , \s_mux1_signals[4][16][26] , 
        \s_mux1_signals[4][16][25] , \s_mux1_signals[4][16][24] , 
        \s_mux1_signals[4][16][23] , \s_mux1_signals[4][16][22] , 
        \s_mux1_signals[4][16][21] , \s_mux1_signals[4][16][20] , 
        \s_mux1_signals[4][16][19] , \s_mux1_signals[4][16][18] , 
        \s_mux1_signals[4][16][17] , \s_mux1_signals[4][16][16] , 
        \s_mux1_signals[4][16][15] , \s_mux1_signals[4][16][14] , 
        \s_mux1_signals[4][16][13] , \s_mux1_signals[4][16][12] , 
        \s_mux1_signals[4][16][11] , \s_mux1_signals[4][16][10] , 
        \s_mux1_signals[4][16][9] , \s_mux1_signals[4][16][8] , 
        \s_mux1_signals[4][16][7] , \s_mux1_signals[4][16][6] , 
        \s_mux1_signals[4][16][5] , \s_mux1_signals[4][16][4] , 
        \s_mux1_signals[4][16][3] , \s_mux1_signals[4][16][2] , 
        \s_mux1_signals[4][16][1] , \s_mux1_signals[4][16][0] }) );
  Mux_NBit_2x1_NBIT_IN32_49 MUX1_4_0 ( .port0({\s_mux1_signals[4][0][31] , 
        \s_mux1_signals[4][0][30] , \s_mux1_signals[4][0][29] , 
        \s_mux1_signals[4][0][28] , \s_mux1_signals[4][0][27] , 
        \s_mux1_signals[4][0][26] , \s_mux1_signals[4][0][25] , 
        \s_mux1_signals[4][0][24] , \s_mux1_signals[4][0][23] , 
        \s_mux1_signals[4][0][22] , \s_mux1_signals[4][0][21] , 
        \s_mux1_signals[4][0][20] , \s_mux1_signals[4][0][19] , 
        \s_mux1_signals[4][0][18] , \s_mux1_signals[4][0][17] , 
        \s_mux1_signals[4][0][16] , \s_mux1_signals[4][0][15] , 
        \s_mux1_signals[4][0][14] , \s_mux1_signals[4][0][13] , 
        \s_mux1_signals[4][0][12] , \s_mux1_signals[4][0][11] , 
        \s_mux1_signals[4][0][10] , \s_mux1_signals[4][0][9] , 
        \s_mux1_signals[4][0][8] , \s_mux1_signals[4][0][7] , 
        \s_mux1_signals[4][0][6] , \s_mux1_signals[4][0][5] , 
        \s_mux1_signals[4][0][4] , \s_mux1_signals[4][0][3] , 
        \s_mux1_signals[4][0][2] , \s_mux1_signals[4][0][1] , 
        \s_mux1_signals[4][0][0] }), .port1({\s_mux1_signals[4][16][31] , 
        \s_mux1_signals[4][16][30] , \s_mux1_signals[4][16][29] , 
        \s_mux1_signals[4][16][28] , \s_mux1_signals[4][16][27] , 
        \s_mux1_signals[4][16][26] , \s_mux1_signals[4][16][25] , 
        \s_mux1_signals[4][16][24] , \s_mux1_signals[4][16][23] , 
        \s_mux1_signals[4][16][22] , \s_mux1_signals[4][16][21] , 
        \s_mux1_signals[4][16][20] , \s_mux1_signals[4][16][19] , 
        \s_mux1_signals[4][16][18] , \s_mux1_signals[4][16][17] , 
        \s_mux1_signals[4][16][16] , \s_mux1_signals[4][16][15] , 
        \s_mux1_signals[4][16][14] , \s_mux1_signals[4][16][13] , 
        \s_mux1_signals[4][16][12] , \s_mux1_signals[4][16][11] , 
        \s_mux1_signals[4][16][10] , \s_mux1_signals[4][16][9] , 
        \s_mux1_signals[4][16][8] , \s_mux1_signals[4][16][7] , 
        \s_mux1_signals[4][16][6] , \s_mux1_signals[4][16][5] , 
        \s_mux1_signals[4][16][4] , \s_mux1_signals[4][16][3] , 
        \s_mux1_signals[4][16][2] , \s_mux1_signals[4][16][1] , 
        \s_mux1_signals[4][16][0] }), .sel(s_addrRd1_Fei_Tmux[4]), .portY(
        RF_out1) );
  Mux_NBit_2x1_NBIT_IN32_48 MUX2_0_0 ( .port0({\s_mux2_signals[0][0][31] , 
        \s_mux2_signals[0][0][30] , \s_mux2_signals[0][0][29] , 
        \s_mux2_signals[0][0][28] , \s_mux2_signals[0][0][27] , 
        \s_mux2_signals[0][0][26] , \s_mux2_signals[0][0][25] , 
        \s_mux2_signals[0][0][24] , \s_mux2_signals[0][0][23] , 
        \s_mux2_signals[0][0][22] , \s_mux2_signals[0][0][21] , 
        \s_mux2_signals[0][0][20] , \s_mux2_signals[0][0][19] , 
        \s_mux2_signals[0][0][18] , \s_mux2_signals[0][0][17] , 
        \s_mux2_signals[0][0][16] , \s_mux2_signals[0][0][15] , 
        \s_mux2_signals[0][0][14] , \s_mux2_signals[0][0][13] , 
        \s_mux2_signals[0][0][12] , \s_mux2_signals[0][0][11] , 
        \s_mux2_signals[0][0][10] , \s_mux2_signals[0][0][9] , 
        \s_mux2_signals[0][0][8] , \s_mux2_signals[0][0][7] , 
        \s_mux2_signals[0][0][6] , \s_mux2_signals[0][0][5] , 
        \s_mux2_signals[0][0][4] , \s_mux2_signals[0][0][3] , 
        \s_mux2_signals[0][0][2] , \s_mux2_signals[0][0][1] , 
        \s_mux2_signals[0][0][0] }), .port1({\s_mux2_signals[0][1][31] , 
        \s_mux2_signals[0][1][30] , \s_mux2_signals[0][1][29] , 
        \s_mux2_signals[0][1][28] , \s_mux2_signals[0][1][27] , 
        \s_mux2_signals[0][1][26] , \s_mux2_signals[0][1][25] , 
        \s_mux2_signals[0][1][24] , \s_mux2_signals[0][1][23] , 
        \s_mux2_signals[0][1][22] , \s_mux2_signals[0][1][21] , 
        \s_mux2_signals[0][1][20] , \s_mux2_signals[0][1][19] , 
        \s_mux2_signals[0][1][18] , \s_mux2_signals[0][1][17] , 
        \s_mux2_signals[0][1][16] , \s_mux2_signals[0][1][15] , 
        \s_mux2_signals[0][1][14] , \s_mux2_signals[0][1][13] , 
        \s_mux2_signals[0][1][12] , \s_mux2_signals[0][1][11] , 
        \s_mux2_signals[0][1][10] , \s_mux2_signals[0][1][9] , 
        \s_mux2_signals[0][1][8] , \s_mux2_signals[0][1][7] , 
        \s_mux2_signals[0][1][6] , \s_mux2_signals[0][1][5] , 
        \s_mux2_signals[0][1][4] , \s_mux2_signals[0][1][3] , 
        \s_mux2_signals[0][1][2] , \s_mux2_signals[0][1][1] , 
        \s_mux2_signals[0][1][0] }), .sel(n25), .portY({
        \s_mux2_signals[1][0][31] , \s_mux2_signals[1][0][30] , 
        \s_mux2_signals[1][0][29] , \s_mux2_signals[1][0][28] , 
        \s_mux2_signals[1][0][27] , \s_mux2_signals[1][0][26] , 
        \s_mux2_signals[1][0][25] , \s_mux2_signals[1][0][24] , 
        \s_mux2_signals[1][0][23] , \s_mux2_signals[1][0][22] , 
        \s_mux2_signals[1][0][21] , \s_mux2_signals[1][0][20] , 
        \s_mux2_signals[1][0][19] , \s_mux2_signals[1][0][18] , 
        \s_mux2_signals[1][0][17] , \s_mux2_signals[1][0][16] , 
        \s_mux2_signals[1][0][15] , \s_mux2_signals[1][0][14] , 
        \s_mux2_signals[1][0][13] , \s_mux2_signals[1][0][12] , 
        \s_mux2_signals[1][0][11] , \s_mux2_signals[1][0][10] , 
        \s_mux2_signals[1][0][9] , \s_mux2_signals[1][0][8] , 
        \s_mux2_signals[1][0][7] , \s_mux2_signals[1][0][6] , 
        \s_mux2_signals[1][0][5] , \s_mux2_signals[1][0][4] , 
        \s_mux2_signals[1][0][3] , \s_mux2_signals[1][0][2] , 
        \s_mux2_signals[1][0][1] , \s_mux2_signals[1][0][0] }) );
  Mux_NBit_2x1_NBIT_IN32_47 MUX2_0_2 ( .port0({\s_mux2_signals[0][2][31] , 
        \s_mux2_signals[0][2][30] , \s_mux2_signals[0][2][29] , 
        \s_mux2_signals[0][2][28] , \s_mux2_signals[0][2][27] , 
        \s_mux2_signals[0][2][26] , \s_mux2_signals[0][2][25] , 
        \s_mux2_signals[0][2][24] , \s_mux2_signals[0][2][23] , 
        \s_mux2_signals[0][2][22] , \s_mux2_signals[0][2][21] , 
        \s_mux2_signals[0][2][20] , \s_mux2_signals[0][2][19] , 
        \s_mux2_signals[0][2][18] , \s_mux2_signals[0][2][17] , 
        \s_mux2_signals[0][2][16] , \s_mux2_signals[0][2][15] , 
        \s_mux2_signals[0][2][14] , \s_mux2_signals[0][2][13] , 
        \s_mux2_signals[0][2][12] , \s_mux2_signals[0][2][11] , 
        \s_mux2_signals[0][2][10] , \s_mux2_signals[0][2][9] , 
        \s_mux2_signals[0][2][8] , \s_mux2_signals[0][2][7] , 
        \s_mux2_signals[0][2][6] , \s_mux2_signals[0][2][5] , 
        \s_mux2_signals[0][2][4] , \s_mux2_signals[0][2][3] , 
        \s_mux2_signals[0][2][2] , \s_mux2_signals[0][2][1] , 
        \s_mux2_signals[0][2][0] }), .port1({\s_mux2_signals[0][3][31] , 
        \s_mux2_signals[0][3][30] , \s_mux2_signals[0][3][29] , 
        \s_mux2_signals[0][3][28] , \s_mux2_signals[0][3][27] , 
        \s_mux2_signals[0][3][26] , \s_mux2_signals[0][3][25] , 
        \s_mux2_signals[0][3][24] , \s_mux2_signals[0][3][23] , 
        \s_mux2_signals[0][3][22] , \s_mux2_signals[0][3][21] , 
        \s_mux2_signals[0][3][20] , \s_mux2_signals[0][3][19] , 
        \s_mux2_signals[0][3][18] , \s_mux2_signals[0][3][17] , 
        \s_mux2_signals[0][3][16] , \s_mux2_signals[0][3][15] , 
        \s_mux2_signals[0][3][14] , \s_mux2_signals[0][3][13] , 
        \s_mux2_signals[0][3][12] , \s_mux2_signals[0][3][11] , 
        \s_mux2_signals[0][3][10] , \s_mux2_signals[0][3][9] , 
        \s_mux2_signals[0][3][8] , \s_mux2_signals[0][3][7] , 
        \s_mux2_signals[0][3][6] , \s_mux2_signals[0][3][5] , 
        \s_mux2_signals[0][3][4] , \s_mux2_signals[0][3][3] , 
        \s_mux2_signals[0][3][2] , \s_mux2_signals[0][3][1] , 
        \s_mux2_signals[0][3][0] }), .sel(n25), .portY({
        \s_mux2_signals[1][2][31] , \s_mux2_signals[1][2][30] , 
        \s_mux2_signals[1][2][29] , \s_mux2_signals[1][2][28] , 
        \s_mux2_signals[1][2][27] , \s_mux2_signals[1][2][26] , 
        \s_mux2_signals[1][2][25] , \s_mux2_signals[1][2][24] , 
        \s_mux2_signals[1][2][23] , \s_mux2_signals[1][2][22] , 
        \s_mux2_signals[1][2][21] , \s_mux2_signals[1][2][20] , 
        \s_mux2_signals[1][2][19] , \s_mux2_signals[1][2][18] , 
        \s_mux2_signals[1][2][17] , \s_mux2_signals[1][2][16] , 
        \s_mux2_signals[1][2][15] , \s_mux2_signals[1][2][14] , 
        \s_mux2_signals[1][2][13] , \s_mux2_signals[1][2][12] , 
        \s_mux2_signals[1][2][11] , \s_mux2_signals[1][2][10] , 
        \s_mux2_signals[1][2][9] , \s_mux2_signals[1][2][8] , 
        \s_mux2_signals[1][2][7] , \s_mux2_signals[1][2][6] , 
        \s_mux2_signals[1][2][5] , \s_mux2_signals[1][2][4] , 
        \s_mux2_signals[1][2][3] , \s_mux2_signals[1][2][2] , 
        \s_mux2_signals[1][2][1] , \s_mux2_signals[1][2][0] }) );
  Mux_NBit_2x1_NBIT_IN32_46 MUX2_0_4 ( .port0({\s_mux2_signals[0][4][31] , 
        \s_mux2_signals[0][4][30] , \s_mux2_signals[0][4][29] , 
        \s_mux2_signals[0][4][28] , \s_mux2_signals[0][4][27] , 
        \s_mux2_signals[0][4][26] , \s_mux2_signals[0][4][25] , 
        \s_mux2_signals[0][4][24] , \s_mux2_signals[0][4][23] , 
        \s_mux2_signals[0][4][22] , \s_mux2_signals[0][4][21] , 
        \s_mux2_signals[0][4][20] , \s_mux2_signals[0][4][19] , 
        \s_mux2_signals[0][4][18] , \s_mux2_signals[0][4][17] , 
        \s_mux2_signals[0][4][16] , \s_mux2_signals[0][4][15] , 
        \s_mux2_signals[0][4][14] , \s_mux2_signals[0][4][13] , 
        \s_mux2_signals[0][4][12] , \s_mux2_signals[0][4][11] , 
        \s_mux2_signals[0][4][10] , \s_mux2_signals[0][4][9] , 
        \s_mux2_signals[0][4][8] , \s_mux2_signals[0][4][7] , 
        \s_mux2_signals[0][4][6] , \s_mux2_signals[0][4][5] , 
        \s_mux2_signals[0][4][4] , \s_mux2_signals[0][4][3] , 
        \s_mux2_signals[0][4][2] , \s_mux2_signals[0][4][1] , 
        \s_mux2_signals[0][4][0] }), .port1({\s_mux2_signals[0][5][31] , 
        \s_mux2_signals[0][5][30] , \s_mux2_signals[0][5][29] , 
        \s_mux2_signals[0][5][28] , \s_mux2_signals[0][5][27] , 
        \s_mux2_signals[0][5][26] , \s_mux2_signals[0][5][25] , 
        \s_mux2_signals[0][5][24] , \s_mux2_signals[0][5][23] , 
        \s_mux2_signals[0][5][22] , \s_mux2_signals[0][5][21] , 
        \s_mux2_signals[0][5][20] , \s_mux2_signals[0][5][19] , 
        \s_mux2_signals[0][5][18] , \s_mux2_signals[0][5][17] , 
        \s_mux2_signals[0][5][16] , \s_mux2_signals[0][5][15] , 
        \s_mux2_signals[0][5][14] , \s_mux2_signals[0][5][13] , 
        \s_mux2_signals[0][5][12] , \s_mux2_signals[0][5][11] , 
        \s_mux2_signals[0][5][10] , \s_mux2_signals[0][5][9] , 
        \s_mux2_signals[0][5][8] , \s_mux2_signals[0][5][7] , 
        \s_mux2_signals[0][5][6] , \s_mux2_signals[0][5][5] , 
        \s_mux2_signals[0][5][4] , \s_mux2_signals[0][5][3] , 
        \s_mux2_signals[0][5][2] , \s_mux2_signals[0][5][1] , 
        \s_mux2_signals[0][5][0] }), .sel(n25), .portY({
        \s_mux2_signals[1][4][31] , \s_mux2_signals[1][4][30] , 
        \s_mux2_signals[1][4][29] , \s_mux2_signals[1][4][28] , 
        \s_mux2_signals[1][4][27] , \s_mux2_signals[1][4][26] , 
        \s_mux2_signals[1][4][25] , \s_mux2_signals[1][4][24] , 
        \s_mux2_signals[1][4][23] , \s_mux2_signals[1][4][22] , 
        \s_mux2_signals[1][4][21] , \s_mux2_signals[1][4][20] , 
        \s_mux2_signals[1][4][19] , \s_mux2_signals[1][4][18] , 
        \s_mux2_signals[1][4][17] , \s_mux2_signals[1][4][16] , 
        \s_mux2_signals[1][4][15] , \s_mux2_signals[1][4][14] , 
        \s_mux2_signals[1][4][13] , \s_mux2_signals[1][4][12] , 
        \s_mux2_signals[1][4][11] , \s_mux2_signals[1][4][10] , 
        \s_mux2_signals[1][4][9] , \s_mux2_signals[1][4][8] , 
        \s_mux2_signals[1][4][7] , \s_mux2_signals[1][4][6] , 
        \s_mux2_signals[1][4][5] , \s_mux2_signals[1][4][4] , 
        \s_mux2_signals[1][4][3] , \s_mux2_signals[1][4][2] , 
        \s_mux2_signals[1][4][1] , \s_mux2_signals[1][4][0] }) );
  Mux_NBit_2x1_NBIT_IN32_45 MUX2_0_6 ( .port0({\s_mux2_signals[0][6][31] , 
        \s_mux2_signals[0][6][30] , \s_mux2_signals[0][6][29] , 
        \s_mux2_signals[0][6][28] , \s_mux2_signals[0][6][27] , 
        \s_mux2_signals[0][6][26] , \s_mux2_signals[0][6][25] , 
        \s_mux2_signals[0][6][24] , \s_mux2_signals[0][6][23] , 
        \s_mux2_signals[0][6][22] , \s_mux2_signals[0][6][21] , 
        \s_mux2_signals[0][6][20] , \s_mux2_signals[0][6][19] , 
        \s_mux2_signals[0][6][18] , \s_mux2_signals[0][6][17] , 
        \s_mux2_signals[0][6][16] , \s_mux2_signals[0][6][15] , 
        \s_mux2_signals[0][6][14] , \s_mux2_signals[0][6][13] , 
        \s_mux2_signals[0][6][12] , \s_mux2_signals[0][6][11] , 
        \s_mux2_signals[0][6][10] , \s_mux2_signals[0][6][9] , 
        \s_mux2_signals[0][6][8] , \s_mux2_signals[0][6][7] , 
        \s_mux2_signals[0][6][6] , \s_mux2_signals[0][6][5] , 
        \s_mux2_signals[0][6][4] , \s_mux2_signals[0][6][3] , 
        \s_mux2_signals[0][6][2] , \s_mux2_signals[0][6][1] , 
        \s_mux2_signals[0][6][0] }), .port1({\s_mux2_signals[0][7][31] , 
        \s_mux2_signals[0][7][30] , \s_mux2_signals[0][7][29] , 
        \s_mux2_signals[0][7][28] , \s_mux2_signals[0][7][27] , 
        \s_mux2_signals[0][7][26] , \s_mux2_signals[0][7][25] , 
        \s_mux2_signals[0][7][24] , \s_mux2_signals[0][7][23] , 
        \s_mux2_signals[0][7][22] , \s_mux2_signals[0][7][21] , 
        \s_mux2_signals[0][7][20] , \s_mux2_signals[0][7][19] , 
        \s_mux2_signals[0][7][18] , \s_mux2_signals[0][7][17] , 
        \s_mux2_signals[0][7][16] , \s_mux2_signals[0][7][15] , 
        \s_mux2_signals[0][7][14] , \s_mux2_signals[0][7][13] , 
        \s_mux2_signals[0][7][12] , \s_mux2_signals[0][7][11] , 
        \s_mux2_signals[0][7][10] , \s_mux2_signals[0][7][9] , 
        \s_mux2_signals[0][7][8] , \s_mux2_signals[0][7][7] , 
        \s_mux2_signals[0][7][6] , \s_mux2_signals[0][7][5] , 
        \s_mux2_signals[0][7][4] , \s_mux2_signals[0][7][3] , 
        \s_mux2_signals[0][7][2] , \s_mux2_signals[0][7][1] , 
        \s_mux2_signals[0][7][0] }), .sel(n25), .portY({
        \s_mux2_signals[1][6][31] , \s_mux2_signals[1][6][30] , 
        \s_mux2_signals[1][6][29] , \s_mux2_signals[1][6][28] , 
        \s_mux2_signals[1][6][27] , \s_mux2_signals[1][6][26] , 
        \s_mux2_signals[1][6][25] , \s_mux2_signals[1][6][24] , 
        \s_mux2_signals[1][6][23] , \s_mux2_signals[1][6][22] , 
        \s_mux2_signals[1][6][21] , \s_mux2_signals[1][6][20] , 
        \s_mux2_signals[1][6][19] , \s_mux2_signals[1][6][18] , 
        \s_mux2_signals[1][6][17] , \s_mux2_signals[1][6][16] , 
        \s_mux2_signals[1][6][15] , \s_mux2_signals[1][6][14] , 
        \s_mux2_signals[1][6][13] , \s_mux2_signals[1][6][12] , 
        \s_mux2_signals[1][6][11] , \s_mux2_signals[1][6][10] , 
        \s_mux2_signals[1][6][9] , \s_mux2_signals[1][6][8] , 
        \s_mux2_signals[1][6][7] , \s_mux2_signals[1][6][6] , 
        \s_mux2_signals[1][6][5] , \s_mux2_signals[1][6][4] , 
        \s_mux2_signals[1][6][3] , \s_mux2_signals[1][6][2] , 
        \s_mux2_signals[1][6][1] , \s_mux2_signals[1][6][0] }) );
  Mux_NBit_2x1_NBIT_IN32_44 MUX2_0_8 ( .port0({\s_mux2_signals[0][8][31] , 
        \s_mux2_signals[0][8][30] , \s_mux2_signals[0][8][29] , 
        \s_mux2_signals[0][8][28] , \s_mux2_signals[0][8][27] , 
        \s_mux2_signals[0][8][26] , \s_mux2_signals[0][8][25] , 
        \s_mux2_signals[0][8][24] , \s_mux2_signals[0][8][23] , 
        \s_mux2_signals[0][8][22] , \s_mux2_signals[0][8][21] , 
        \s_mux2_signals[0][8][20] , \s_mux2_signals[0][8][19] , 
        \s_mux2_signals[0][8][18] , \s_mux2_signals[0][8][17] , 
        \s_mux2_signals[0][8][16] , \s_mux2_signals[0][8][15] , 
        \s_mux2_signals[0][8][14] , \s_mux2_signals[0][8][13] , 
        \s_mux2_signals[0][8][12] , \s_mux2_signals[0][8][11] , 
        \s_mux2_signals[0][8][10] , \s_mux2_signals[0][8][9] , 
        \s_mux2_signals[0][8][8] , \s_mux2_signals[0][8][7] , 
        \s_mux2_signals[0][8][6] , \s_mux2_signals[0][8][5] , 
        \s_mux2_signals[0][8][4] , \s_mux2_signals[0][8][3] , 
        \s_mux2_signals[0][8][2] , \s_mux2_signals[0][8][1] , 
        \s_mux2_signals[0][8][0] }), .port1({\s_mux2_signals[0][9][31] , 
        \s_mux2_signals[0][9][30] , \s_mux2_signals[0][9][29] , 
        \s_mux2_signals[0][9][28] , \s_mux2_signals[0][9][27] , 
        \s_mux2_signals[0][9][26] , \s_mux2_signals[0][9][25] , 
        \s_mux2_signals[0][9][24] , \s_mux2_signals[0][9][23] , 
        \s_mux2_signals[0][9][22] , \s_mux2_signals[0][9][21] , 
        \s_mux2_signals[0][9][20] , \s_mux2_signals[0][9][19] , 
        \s_mux2_signals[0][9][18] , \s_mux2_signals[0][9][17] , 
        \s_mux2_signals[0][9][16] , \s_mux2_signals[0][9][15] , 
        \s_mux2_signals[0][9][14] , \s_mux2_signals[0][9][13] , 
        \s_mux2_signals[0][9][12] , \s_mux2_signals[0][9][11] , 
        \s_mux2_signals[0][9][10] , \s_mux2_signals[0][9][9] , 
        \s_mux2_signals[0][9][8] , \s_mux2_signals[0][9][7] , 
        \s_mux2_signals[0][9][6] , \s_mux2_signals[0][9][5] , 
        \s_mux2_signals[0][9][4] , \s_mux2_signals[0][9][3] , 
        \s_mux2_signals[0][9][2] , \s_mux2_signals[0][9][1] , 
        \s_mux2_signals[0][9][0] }), .sel(n25), .portY({
        \s_mux2_signals[1][8][31] , \s_mux2_signals[1][8][30] , 
        \s_mux2_signals[1][8][29] , \s_mux2_signals[1][8][28] , 
        \s_mux2_signals[1][8][27] , \s_mux2_signals[1][8][26] , 
        \s_mux2_signals[1][8][25] , \s_mux2_signals[1][8][24] , 
        \s_mux2_signals[1][8][23] , \s_mux2_signals[1][8][22] , 
        \s_mux2_signals[1][8][21] , \s_mux2_signals[1][8][20] , 
        \s_mux2_signals[1][8][19] , \s_mux2_signals[1][8][18] , 
        \s_mux2_signals[1][8][17] , \s_mux2_signals[1][8][16] , 
        \s_mux2_signals[1][8][15] , \s_mux2_signals[1][8][14] , 
        \s_mux2_signals[1][8][13] , \s_mux2_signals[1][8][12] , 
        \s_mux2_signals[1][8][11] , \s_mux2_signals[1][8][10] , 
        \s_mux2_signals[1][8][9] , \s_mux2_signals[1][8][8] , 
        \s_mux2_signals[1][8][7] , \s_mux2_signals[1][8][6] , 
        \s_mux2_signals[1][8][5] , \s_mux2_signals[1][8][4] , 
        \s_mux2_signals[1][8][3] , \s_mux2_signals[1][8][2] , 
        \s_mux2_signals[1][8][1] , \s_mux2_signals[1][8][0] }) );
  Mux_NBit_2x1_NBIT_IN32_43 MUX2_0_10 ( .port0({\s_mux2_signals[0][10][31] , 
        \s_mux2_signals[0][10][30] , \s_mux2_signals[0][10][29] , 
        \s_mux2_signals[0][10][28] , \s_mux2_signals[0][10][27] , 
        \s_mux2_signals[0][10][26] , \s_mux2_signals[0][10][25] , 
        \s_mux2_signals[0][10][24] , \s_mux2_signals[0][10][23] , 
        \s_mux2_signals[0][10][22] , \s_mux2_signals[0][10][21] , 
        \s_mux2_signals[0][10][20] , \s_mux2_signals[0][10][19] , 
        \s_mux2_signals[0][10][18] , \s_mux2_signals[0][10][17] , 
        \s_mux2_signals[0][10][16] , \s_mux2_signals[0][10][15] , 
        \s_mux2_signals[0][10][14] , \s_mux2_signals[0][10][13] , 
        \s_mux2_signals[0][10][12] , \s_mux2_signals[0][10][11] , 
        \s_mux2_signals[0][10][10] , \s_mux2_signals[0][10][9] , 
        \s_mux2_signals[0][10][8] , \s_mux2_signals[0][10][7] , 
        \s_mux2_signals[0][10][6] , \s_mux2_signals[0][10][5] , 
        \s_mux2_signals[0][10][4] , \s_mux2_signals[0][10][3] , 
        \s_mux2_signals[0][10][2] , \s_mux2_signals[0][10][1] , 
        \s_mux2_signals[0][10][0] }), .port1({\s_mux2_signals[0][11][31] , 
        \s_mux2_signals[0][11][30] , \s_mux2_signals[0][11][29] , 
        \s_mux2_signals[0][11][28] , \s_mux2_signals[0][11][27] , 
        \s_mux2_signals[0][11][26] , \s_mux2_signals[0][11][25] , 
        \s_mux2_signals[0][11][24] , \s_mux2_signals[0][11][23] , 
        \s_mux2_signals[0][11][22] , \s_mux2_signals[0][11][21] , 
        \s_mux2_signals[0][11][20] , \s_mux2_signals[0][11][19] , 
        \s_mux2_signals[0][11][18] , \s_mux2_signals[0][11][17] , 
        \s_mux2_signals[0][11][16] , \s_mux2_signals[0][11][15] , 
        \s_mux2_signals[0][11][14] , \s_mux2_signals[0][11][13] , 
        \s_mux2_signals[0][11][12] , \s_mux2_signals[0][11][11] , 
        \s_mux2_signals[0][11][10] , \s_mux2_signals[0][11][9] , 
        \s_mux2_signals[0][11][8] , \s_mux2_signals[0][11][7] , 
        \s_mux2_signals[0][11][6] , \s_mux2_signals[0][11][5] , 
        \s_mux2_signals[0][11][4] , \s_mux2_signals[0][11][3] , 
        \s_mux2_signals[0][11][2] , \s_mux2_signals[0][11][1] , 
        \s_mux2_signals[0][11][0] }), .sel(n25), .portY({
        \s_mux2_signals[1][10][31] , \s_mux2_signals[1][10][30] , 
        \s_mux2_signals[1][10][29] , \s_mux2_signals[1][10][28] , 
        \s_mux2_signals[1][10][27] , \s_mux2_signals[1][10][26] , 
        \s_mux2_signals[1][10][25] , \s_mux2_signals[1][10][24] , 
        \s_mux2_signals[1][10][23] , \s_mux2_signals[1][10][22] , 
        \s_mux2_signals[1][10][21] , \s_mux2_signals[1][10][20] , 
        \s_mux2_signals[1][10][19] , \s_mux2_signals[1][10][18] , 
        \s_mux2_signals[1][10][17] , \s_mux2_signals[1][10][16] , 
        \s_mux2_signals[1][10][15] , \s_mux2_signals[1][10][14] , 
        \s_mux2_signals[1][10][13] , \s_mux2_signals[1][10][12] , 
        \s_mux2_signals[1][10][11] , \s_mux2_signals[1][10][10] , 
        \s_mux2_signals[1][10][9] , \s_mux2_signals[1][10][8] , 
        \s_mux2_signals[1][10][7] , \s_mux2_signals[1][10][6] , 
        \s_mux2_signals[1][10][5] , \s_mux2_signals[1][10][4] , 
        \s_mux2_signals[1][10][3] , \s_mux2_signals[1][10][2] , 
        \s_mux2_signals[1][10][1] , \s_mux2_signals[1][10][0] }) );
  Mux_NBit_2x1_NBIT_IN32_42 MUX2_0_12 ( .port0({\s_mux2_signals[0][12][31] , 
        \s_mux2_signals[0][12][30] , \s_mux2_signals[0][12][29] , 
        \s_mux2_signals[0][12][28] , \s_mux2_signals[0][12][27] , 
        \s_mux2_signals[0][12][26] , \s_mux2_signals[0][12][25] , 
        \s_mux2_signals[0][12][24] , \s_mux2_signals[0][12][23] , 
        \s_mux2_signals[0][12][22] , \s_mux2_signals[0][12][21] , 
        \s_mux2_signals[0][12][20] , \s_mux2_signals[0][12][19] , 
        \s_mux2_signals[0][12][18] , \s_mux2_signals[0][12][17] , 
        \s_mux2_signals[0][12][16] , \s_mux2_signals[0][12][15] , 
        \s_mux2_signals[0][12][14] , \s_mux2_signals[0][12][13] , 
        \s_mux2_signals[0][12][12] , \s_mux2_signals[0][12][11] , 
        \s_mux2_signals[0][12][10] , \s_mux2_signals[0][12][9] , 
        \s_mux2_signals[0][12][8] , \s_mux2_signals[0][12][7] , 
        \s_mux2_signals[0][12][6] , \s_mux2_signals[0][12][5] , 
        \s_mux2_signals[0][12][4] , \s_mux2_signals[0][12][3] , 
        \s_mux2_signals[0][12][2] , \s_mux2_signals[0][12][1] , 
        \s_mux2_signals[0][12][0] }), .port1({\s_mux2_signals[0][13][31] , 
        \s_mux2_signals[0][13][30] , \s_mux2_signals[0][13][29] , 
        \s_mux2_signals[0][13][28] , \s_mux2_signals[0][13][27] , 
        \s_mux2_signals[0][13][26] , \s_mux2_signals[0][13][25] , 
        \s_mux2_signals[0][13][24] , \s_mux2_signals[0][13][23] , 
        \s_mux2_signals[0][13][22] , \s_mux2_signals[0][13][21] , 
        \s_mux2_signals[0][13][20] , \s_mux2_signals[0][13][19] , 
        \s_mux2_signals[0][13][18] , \s_mux2_signals[0][13][17] , 
        \s_mux2_signals[0][13][16] , \s_mux2_signals[0][13][15] , 
        \s_mux2_signals[0][13][14] , \s_mux2_signals[0][13][13] , 
        \s_mux2_signals[0][13][12] , \s_mux2_signals[0][13][11] , 
        \s_mux2_signals[0][13][10] , \s_mux2_signals[0][13][9] , 
        \s_mux2_signals[0][13][8] , \s_mux2_signals[0][13][7] , 
        \s_mux2_signals[0][13][6] , \s_mux2_signals[0][13][5] , 
        \s_mux2_signals[0][13][4] , \s_mux2_signals[0][13][3] , 
        \s_mux2_signals[0][13][2] , \s_mux2_signals[0][13][1] , 
        \s_mux2_signals[0][13][0] }), .sel(n25), .portY({
        \s_mux2_signals[1][12][31] , \s_mux2_signals[1][12][30] , 
        \s_mux2_signals[1][12][29] , \s_mux2_signals[1][12][28] , 
        \s_mux2_signals[1][12][27] , \s_mux2_signals[1][12][26] , 
        \s_mux2_signals[1][12][25] , \s_mux2_signals[1][12][24] , 
        \s_mux2_signals[1][12][23] , \s_mux2_signals[1][12][22] , 
        \s_mux2_signals[1][12][21] , \s_mux2_signals[1][12][20] , 
        \s_mux2_signals[1][12][19] , \s_mux2_signals[1][12][18] , 
        \s_mux2_signals[1][12][17] , \s_mux2_signals[1][12][16] , 
        \s_mux2_signals[1][12][15] , \s_mux2_signals[1][12][14] , 
        \s_mux2_signals[1][12][13] , \s_mux2_signals[1][12][12] , 
        \s_mux2_signals[1][12][11] , \s_mux2_signals[1][12][10] , 
        \s_mux2_signals[1][12][9] , \s_mux2_signals[1][12][8] , 
        \s_mux2_signals[1][12][7] , \s_mux2_signals[1][12][6] , 
        \s_mux2_signals[1][12][5] , \s_mux2_signals[1][12][4] , 
        \s_mux2_signals[1][12][3] , \s_mux2_signals[1][12][2] , 
        \s_mux2_signals[1][12][1] , \s_mux2_signals[1][12][0] }) );
  Mux_NBit_2x1_NBIT_IN32_41 MUX2_0_14 ( .port0({\s_mux2_signals[0][14][31] , 
        \s_mux2_signals[0][14][30] , \s_mux2_signals[0][14][29] , 
        \s_mux2_signals[0][14][28] , \s_mux2_signals[0][14][27] , 
        \s_mux2_signals[0][14][26] , \s_mux2_signals[0][14][25] , 
        \s_mux2_signals[0][14][24] , \s_mux2_signals[0][14][23] , 
        \s_mux2_signals[0][14][22] , \s_mux2_signals[0][14][21] , 
        \s_mux2_signals[0][14][20] , \s_mux2_signals[0][14][19] , 
        \s_mux2_signals[0][14][18] , \s_mux2_signals[0][14][17] , 
        \s_mux2_signals[0][14][16] , \s_mux2_signals[0][14][15] , 
        \s_mux2_signals[0][14][14] , \s_mux2_signals[0][14][13] , 
        \s_mux2_signals[0][14][12] , \s_mux2_signals[0][14][11] , 
        \s_mux2_signals[0][14][10] , \s_mux2_signals[0][14][9] , 
        \s_mux2_signals[0][14][8] , \s_mux2_signals[0][14][7] , 
        \s_mux2_signals[0][14][6] , \s_mux2_signals[0][14][5] , 
        \s_mux2_signals[0][14][4] , \s_mux2_signals[0][14][3] , 
        \s_mux2_signals[0][14][2] , \s_mux2_signals[0][14][1] , 
        \s_mux2_signals[0][14][0] }), .port1({\s_mux2_signals[0][15][31] , 
        \s_mux2_signals[0][15][30] , \s_mux2_signals[0][15][29] , 
        \s_mux2_signals[0][15][28] , \s_mux2_signals[0][15][27] , 
        \s_mux2_signals[0][15][26] , \s_mux2_signals[0][15][25] , 
        \s_mux2_signals[0][15][24] , \s_mux2_signals[0][15][23] , 
        \s_mux2_signals[0][15][22] , \s_mux2_signals[0][15][21] , 
        \s_mux2_signals[0][15][20] , \s_mux2_signals[0][15][19] , 
        \s_mux2_signals[0][15][18] , \s_mux2_signals[0][15][17] , 
        \s_mux2_signals[0][15][16] , \s_mux2_signals[0][15][15] , 
        \s_mux2_signals[0][15][14] , \s_mux2_signals[0][15][13] , 
        \s_mux2_signals[0][15][12] , \s_mux2_signals[0][15][11] , 
        \s_mux2_signals[0][15][10] , \s_mux2_signals[0][15][9] , 
        \s_mux2_signals[0][15][8] , \s_mux2_signals[0][15][7] , 
        \s_mux2_signals[0][15][6] , \s_mux2_signals[0][15][5] , 
        \s_mux2_signals[0][15][4] , \s_mux2_signals[0][15][3] , 
        \s_mux2_signals[0][15][2] , \s_mux2_signals[0][15][1] , 
        \s_mux2_signals[0][15][0] }), .sel(n26), .portY({
        \s_mux2_signals[1][14][31] , \s_mux2_signals[1][14][30] , 
        \s_mux2_signals[1][14][29] , \s_mux2_signals[1][14][28] , 
        \s_mux2_signals[1][14][27] , \s_mux2_signals[1][14][26] , 
        \s_mux2_signals[1][14][25] , \s_mux2_signals[1][14][24] , 
        \s_mux2_signals[1][14][23] , \s_mux2_signals[1][14][22] , 
        \s_mux2_signals[1][14][21] , \s_mux2_signals[1][14][20] , 
        \s_mux2_signals[1][14][19] , \s_mux2_signals[1][14][18] , 
        \s_mux2_signals[1][14][17] , \s_mux2_signals[1][14][16] , 
        \s_mux2_signals[1][14][15] , \s_mux2_signals[1][14][14] , 
        \s_mux2_signals[1][14][13] , \s_mux2_signals[1][14][12] , 
        \s_mux2_signals[1][14][11] , \s_mux2_signals[1][14][10] , 
        \s_mux2_signals[1][14][9] , \s_mux2_signals[1][14][8] , 
        \s_mux2_signals[1][14][7] , \s_mux2_signals[1][14][6] , 
        \s_mux2_signals[1][14][5] , \s_mux2_signals[1][14][4] , 
        \s_mux2_signals[1][14][3] , \s_mux2_signals[1][14][2] , 
        \s_mux2_signals[1][14][1] , \s_mux2_signals[1][14][0] }) );
  Mux_NBit_2x1_NBIT_IN32_40 MUX2_0_16 ( .port0({\s_mux2_signals[0][16][31] , 
        \s_mux2_signals[0][16][30] , \s_mux2_signals[0][16][29] , 
        \s_mux2_signals[0][16][28] , \s_mux2_signals[0][16][27] , 
        \s_mux2_signals[0][16][26] , \s_mux2_signals[0][16][25] , 
        \s_mux2_signals[0][16][24] , \s_mux2_signals[0][16][23] , 
        \s_mux2_signals[0][16][22] , \s_mux2_signals[0][16][21] , 
        \s_mux2_signals[0][16][20] , \s_mux2_signals[0][16][19] , 
        \s_mux2_signals[0][16][18] , \s_mux2_signals[0][16][17] , 
        \s_mux2_signals[0][16][16] , \s_mux2_signals[0][16][15] , 
        \s_mux2_signals[0][16][14] , \s_mux2_signals[0][16][13] , 
        \s_mux2_signals[0][16][12] , \s_mux2_signals[0][16][11] , 
        \s_mux2_signals[0][16][10] , \s_mux2_signals[0][16][9] , 
        \s_mux2_signals[0][16][8] , \s_mux2_signals[0][16][7] , 
        \s_mux2_signals[0][16][6] , \s_mux2_signals[0][16][5] , 
        \s_mux2_signals[0][16][4] , \s_mux2_signals[0][16][3] , 
        \s_mux2_signals[0][16][2] , \s_mux2_signals[0][16][1] , 
        \s_mux2_signals[0][16][0] }), .port1({\s_mux2_signals[0][17][31] , 
        \s_mux2_signals[0][17][30] , \s_mux2_signals[0][17][29] , 
        \s_mux2_signals[0][17][28] , \s_mux2_signals[0][17][27] , 
        \s_mux2_signals[0][17][26] , \s_mux2_signals[0][17][25] , 
        \s_mux2_signals[0][17][24] , \s_mux2_signals[0][17][23] , 
        \s_mux2_signals[0][17][22] , \s_mux2_signals[0][17][21] , 
        \s_mux2_signals[0][17][20] , \s_mux2_signals[0][17][19] , 
        \s_mux2_signals[0][17][18] , \s_mux2_signals[0][17][17] , 
        \s_mux2_signals[0][17][16] , \s_mux2_signals[0][17][15] , 
        \s_mux2_signals[0][17][14] , \s_mux2_signals[0][17][13] , 
        \s_mux2_signals[0][17][12] , \s_mux2_signals[0][17][11] , 
        \s_mux2_signals[0][17][10] , \s_mux2_signals[0][17][9] , 
        \s_mux2_signals[0][17][8] , \s_mux2_signals[0][17][7] , 
        \s_mux2_signals[0][17][6] , \s_mux2_signals[0][17][5] , 
        \s_mux2_signals[0][17][4] , \s_mux2_signals[0][17][3] , 
        \s_mux2_signals[0][17][2] , \s_mux2_signals[0][17][1] , 
        \s_mux2_signals[0][17][0] }), .sel(n26), .portY({
        \s_mux2_signals[1][16][31] , \s_mux2_signals[1][16][30] , 
        \s_mux2_signals[1][16][29] , \s_mux2_signals[1][16][28] , 
        \s_mux2_signals[1][16][27] , \s_mux2_signals[1][16][26] , 
        \s_mux2_signals[1][16][25] , \s_mux2_signals[1][16][24] , 
        \s_mux2_signals[1][16][23] , \s_mux2_signals[1][16][22] , 
        \s_mux2_signals[1][16][21] , \s_mux2_signals[1][16][20] , 
        \s_mux2_signals[1][16][19] , \s_mux2_signals[1][16][18] , 
        \s_mux2_signals[1][16][17] , \s_mux2_signals[1][16][16] , 
        \s_mux2_signals[1][16][15] , \s_mux2_signals[1][16][14] , 
        \s_mux2_signals[1][16][13] , \s_mux2_signals[1][16][12] , 
        \s_mux2_signals[1][16][11] , \s_mux2_signals[1][16][10] , 
        \s_mux2_signals[1][16][9] , \s_mux2_signals[1][16][8] , 
        \s_mux2_signals[1][16][7] , \s_mux2_signals[1][16][6] , 
        \s_mux2_signals[1][16][5] , \s_mux2_signals[1][16][4] , 
        \s_mux2_signals[1][16][3] , \s_mux2_signals[1][16][2] , 
        \s_mux2_signals[1][16][1] , \s_mux2_signals[1][16][0] }) );
  Mux_NBit_2x1_NBIT_IN32_39 MUX2_0_18 ( .port0({\s_mux2_signals[0][18][31] , 
        \s_mux2_signals[0][18][30] , \s_mux2_signals[0][18][29] , 
        \s_mux2_signals[0][18][28] , \s_mux2_signals[0][18][27] , 
        \s_mux2_signals[0][18][26] , \s_mux2_signals[0][18][25] , 
        \s_mux2_signals[0][18][24] , \s_mux2_signals[0][18][23] , 
        \s_mux2_signals[0][18][22] , \s_mux2_signals[0][18][21] , 
        \s_mux2_signals[0][18][20] , \s_mux2_signals[0][18][19] , 
        \s_mux2_signals[0][18][18] , \s_mux2_signals[0][18][17] , 
        \s_mux2_signals[0][18][16] , \s_mux2_signals[0][18][15] , 
        \s_mux2_signals[0][18][14] , \s_mux2_signals[0][18][13] , 
        \s_mux2_signals[0][18][12] , \s_mux2_signals[0][18][11] , 
        \s_mux2_signals[0][18][10] , \s_mux2_signals[0][18][9] , 
        \s_mux2_signals[0][18][8] , \s_mux2_signals[0][18][7] , 
        \s_mux2_signals[0][18][6] , \s_mux2_signals[0][18][5] , 
        \s_mux2_signals[0][18][4] , \s_mux2_signals[0][18][3] , 
        \s_mux2_signals[0][18][2] , \s_mux2_signals[0][18][1] , 
        \s_mux2_signals[0][18][0] }), .port1({\s_mux2_signals[0][19][31] , 
        \s_mux2_signals[0][19][30] , \s_mux2_signals[0][19][29] , 
        \s_mux2_signals[0][19][28] , \s_mux2_signals[0][19][27] , 
        \s_mux2_signals[0][19][26] , \s_mux2_signals[0][19][25] , 
        \s_mux2_signals[0][19][24] , \s_mux2_signals[0][19][23] , 
        \s_mux2_signals[0][19][22] , \s_mux2_signals[0][19][21] , 
        \s_mux2_signals[0][19][20] , \s_mux2_signals[0][19][19] , 
        \s_mux2_signals[0][19][18] , \s_mux2_signals[0][19][17] , 
        \s_mux2_signals[0][19][16] , \s_mux2_signals[0][19][15] , 
        \s_mux2_signals[0][19][14] , \s_mux2_signals[0][19][13] , 
        \s_mux2_signals[0][19][12] , \s_mux2_signals[0][19][11] , 
        \s_mux2_signals[0][19][10] , \s_mux2_signals[0][19][9] , 
        \s_mux2_signals[0][19][8] , \s_mux2_signals[0][19][7] , 
        \s_mux2_signals[0][19][6] , \s_mux2_signals[0][19][5] , 
        \s_mux2_signals[0][19][4] , \s_mux2_signals[0][19][3] , 
        \s_mux2_signals[0][19][2] , \s_mux2_signals[0][19][1] , 
        \s_mux2_signals[0][19][0] }), .sel(n26), .portY({
        \s_mux2_signals[1][18][31] , \s_mux2_signals[1][18][30] , 
        \s_mux2_signals[1][18][29] , \s_mux2_signals[1][18][28] , 
        \s_mux2_signals[1][18][27] , \s_mux2_signals[1][18][26] , 
        \s_mux2_signals[1][18][25] , \s_mux2_signals[1][18][24] , 
        \s_mux2_signals[1][18][23] , \s_mux2_signals[1][18][22] , 
        \s_mux2_signals[1][18][21] , \s_mux2_signals[1][18][20] , 
        \s_mux2_signals[1][18][19] , \s_mux2_signals[1][18][18] , 
        \s_mux2_signals[1][18][17] , \s_mux2_signals[1][18][16] , 
        \s_mux2_signals[1][18][15] , \s_mux2_signals[1][18][14] , 
        \s_mux2_signals[1][18][13] , \s_mux2_signals[1][18][12] , 
        \s_mux2_signals[1][18][11] , \s_mux2_signals[1][18][10] , 
        \s_mux2_signals[1][18][9] , \s_mux2_signals[1][18][8] , 
        \s_mux2_signals[1][18][7] , \s_mux2_signals[1][18][6] , 
        \s_mux2_signals[1][18][5] , \s_mux2_signals[1][18][4] , 
        \s_mux2_signals[1][18][3] , \s_mux2_signals[1][18][2] , 
        \s_mux2_signals[1][18][1] , \s_mux2_signals[1][18][0] }) );
  Mux_NBit_2x1_NBIT_IN32_38 MUX2_0_20 ( .port0({\s_mux2_signals[0][20][31] , 
        \s_mux2_signals[0][20][30] , \s_mux2_signals[0][20][29] , 
        \s_mux2_signals[0][20][28] , \s_mux2_signals[0][20][27] , 
        \s_mux2_signals[0][20][26] , \s_mux2_signals[0][20][25] , 
        \s_mux2_signals[0][20][24] , \s_mux2_signals[0][20][23] , 
        \s_mux2_signals[0][20][22] , \s_mux2_signals[0][20][21] , 
        \s_mux2_signals[0][20][20] , \s_mux2_signals[0][20][19] , 
        \s_mux2_signals[0][20][18] , \s_mux2_signals[0][20][17] , 
        \s_mux2_signals[0][20][16] , \s_mux2_signals[0][20][15] , 
        \s_mux2_signals[0][20][14] , \s_mux2_signals[0][20][13] , 
        \s_mux2_signals[0][20][12] , \s_mux2_signals[0][20][11] , 
        \s_mux2_signals[0][20][10] , \s_mux2_signals[0][20][9] , 
        \s_mux2_signals[0][20][8] , \s_mux2_signals[0][20][7] , 
        \s_mux2_signals[0][20][6] , \s_mux2_signals[0][20][5] , 
        \s_mux2_signals[0][20][4] , \s_mux2_signals[0][20][3] , 
        \s_mux2_signals[0][20][2] , \s_mux2_signals[0][20][1] , 
        \s_mux2_signals[0][20][0] }), .port1({\s_mux2_signals[0][21][31] , 
        \s_mux2_signals[0][21][30] , \s_mux2_signals[0][21][29] , 
        \s_mux2_signals[0][21][28] , \s_mux2_signals[0][21][27] , 
        \s_mux2_signals[0][21][26] , \s_mux2_signals[0][21][25] , 
        \s_mux2_signals[0][21][24] , \s_mux2_signals[0][21][23] , 
        \s_mux2_signals[0][21][22] , \s_mux2_signals[0][21][21] , 
        \s_mux2_signals[0][21][20] , \s_mux2_signals[0][21][19] , 
        \s_mux2_signals[0][21][18] , \s_mux2_signals[0][21][17] , 
        \s_mux2_signals[0][21][16] , \s_mux2_signals[0][21][15] , 
        \s_mux2_signals[0][21][14] , \s_mux2_signals[0][21][13] , 
        \s_mux2_signals[0][21][12] , \s_mux2_signals[0][21][11] , 
        \s_mux2_signals[0][21][10] , \s_mux2_signals[0][21][9] , 
        \s_mux2_signals[0][21][8] , \s_mux2_signals[0][21][7] , 
        \s_mux2_signals[0][21][6] , \s_mux2_signals[0][21][5] , 
        \s_mux2_signals[0][21][4] , \s_mux2_signals[0][21][3] , 
        \s_mux2_signals[0][21][2] , \s_mux2_signals[0][21][1] , 
        \s_mux2_signals[0][21][0] }), .sel(n26), .portY({
        \s_mux2_signals[1][20][31] , \s_mux2_signals[1][20][30] , 
        \s_mux2_signals[1][20][29] , \s_mux2_signals[1][20][28] , 
        \s_mux2_signals[1][20][27] , \s_mux2_signals[1][20][26] , 
        \s_mux2_signals[1][20][25] , \s_mux2_signals[1][20][24] , 
        \s_mux2_signals[1][20][23] , \s_mux2_signals[1][20][22] , 
        \s_mux2_signals[1][20][21] , \s_mux2_signals[1][20][20] , 
        \s_mux2_signals[1][20][19] , \s_mux2_signals[1][20][18] , 
        \s_mux2_signals[1][20][17] , \s_mux2_signals[1][20][16] , 
        \s_mux2_signals[1][20][15] , \s_mux2_signals[1][20][14] , 
        \s_mux2_signals[1][20][13] , \s_mux2_signals[1][20][12] , 
        \s_mux2_signals[1][20][11] , \s_mux2_signals[1][20][10] , 
        \s_mux2_signals[1][20][9] , \s_mux2_signals[1][20][8] , 
        \s_mux2_signals[1][20][7] , \s_mux2_signals[1][20][6] , 
        \s_mux2_signals[1][20][5] , \s_mux2_signals[1][20][4] , 
        \s_mux2_signals[1][20][3] , \s_mux2_signals[1][20][2] , 
        \s_mux2_signals[1][20][1] , \s_mux2_signals[1][20][0] }) );
  Mux_NBit_2x1_NBIT_IN32_37 MUX2_0_22 ( .port0({\s_mux2_signals[0][22][31] , 
        \s_mux2_signals[0][22][30] , \s_mux2_signals[0][22][29] , 
        \s_mux2_signals[0][22][28] , \s_mux2_signals[0][22][27] , 
        \s_mux2_signals[0][22][26] , \s_mux2_signals[0][22][25] , 
        \s_mux2_signals[0][22][24] , \s_mux2_signals[0][22][23] , 
        \s_mux2_signals[0][22][22] , \s_mux2_signals[0][22][21] , 
        \s_mux2_signals[0][22][20] , \s_mux2_signals[0][22][19] , 
        \s_mux2_signals[0][22][18] , \s_mux2_signals[0][22][17] , 
        \s_mux2_signals[0][22][16] , \s_mux2_signals[0][22][15] , 
        \s_mux2_signals[0][22][14] , \s_mux2_signals[0][22][13] , 
        \s_mux2_signals[0][22][12] , \s_mux2_signals[0][22][11] , 
        \s_mux2_signals[0][22][10] , \s_mux2_signals[0][22][9] , 
        \s_mux2_signals[0][22][8] , \s_mux2_signals[0][22][7] , 
        \s_mux2_signals[0][22][6] , \s_mux2_signals[0][22][5] , 
        \s_mux2_signals[0][22][4] , \s_mux2_signals[0][22][3] , 
        \s_mux2_signals[0][22][2] , \s_mux2_signals[0][22][1] , 
        \s_mux2_signals[0][22][0] }), .port1({\s_mux2_signals[0][23][31] , 
        \s_mux2_signals[0][23][30] , \s_mux2_signals[0][23][29] , 
        \s_mux2_signals[0][23][28] , \s_mux2_signals[0][23][27] , 
        \s_mux2_signals[0][23][26] , \s_mux2_signals[0][23][25] , 
        \s_mux2_signals[0][23][24] , \s_mux2_signals[0][23][23] , 
        \s_mux2_signals[0][23][22] , \s_mux2_signals[0][23][21] , 
        \s_mux2_signals[0][23][20] , \s_mux2_signals[0][23][19] , 
        \s_mux2_signals[0][23][18] , \s_mux2_signals[0][23][17] , 
        \s_mux2_signals[0][23][16] , \s_mux2_signals[0][23][15] , 
        \s_mux2_signals[0][23][14] , \s_mux2_signals[0][23][13] , 
        \s_mux2_signals[0][23][12] , \s_mux2_signals[0][23][11] , 
        \s_mux2_signals[0][23][10] , \s_mux2_signals[0][23][9] , 
        \s_mux2_signals[0][23][8] , \s_mux2_signals[0][23][7] , 
        \s_mux2_signals[0][23][6] , \s_mux2_signals[0][23][5] , 
        \s_mux2_signals[0][23][4] , \s_mux2_signals[0][23][3] , 
        \s_mux2_signals[0][23][2] , \s_mux2_signals[0][23][1] , 
        \s_mux2_signals[0][23][0] }), .sel(n26), .portY({
        \s_mux2_signals[1][22][31] , \s_mux2_signals[1][22][30] , 
        \s_mux2_signals[1][22][29] , \s_mux2_signals[1][22][28] , 
        \s_mux2_signals[1][22][27] , \s_mux2_signals[1][22][26] , 
        \s_mux2_signals[1][22][25] , \s_mux2_signals[1][22][24] , 
        \s_mux2_signals[1][22][23] , \s_mux2_signals[1][22][22] , 
        \s_mux2_signals[1][22][21] , \s_mux2_signals[1][22][20] , 
        \s_mux2_signals[1][22][19] , \s_mux2_signals[1][22][18] , 
        \s_mux2_signals[1][22][17] , \s_mux2_signals[1][22][16] , 
        \s_mux2_signals[1][22][15] , \s_mux2_signals[1][22][14] , 
        \s_mux2_signals[1][22][13] , \s_mux2_signals[1][22][12] , 
        \s_mux2_signals[1][22][11] , \s_mux2_signals[1][22][10] , 
        \s_mux2_signals[1][22][9] , \s_mux2_signals[1][22][8] , 
        \s_mux2_signals[1][22][7] , \s_mux2_signals[1][22][6] , 
        \s_mux2_signals[1][22][5] , \s_mux2_signals[1][22][4] , 
        \s_mux2_signals[1][22][3] , \s_mux2_signals[1][22][2] , 
        \s_mux2_signals[1][22][1] , \s_mux2_signals[1][22][0] }) );
  Mux_NBit_2x1_NBIT_IN32_36 MUX2_0_24 ( .port0({\s_mux2_signals[0][24][31] , 
        \s_mux2_signals[0][24][30] , \s_mux2_signals[0][24][29] , 
        \s_mux2_signals[0][24][28] , \s_mux2_signals[0][24][27] , 
        \s_mux2_signals[0][24][26] , \s_mux2_signals[0][24][25] , 
        \s_mux2_signals[0][24][24] , \s_mux2_signals[0][24][23] , 
        \s_mux2_signals[0][24][22] , \s_mux2_signals[0][24][21] , 
        \s_mux2_signals[0][24][20] , \s_mux2_signals[0][24][19] , 
        \s_mux2_signals[0][24][18] , \s_mux2_signals[0][24][17] , 
        \s_mux2_signals[0][24][16] , \s_mux2_signals[0][24][15] , 
        \s_mux2_signals[0][24][14] , \s_mux2_signals[0][24][13] , 
        \s_mux2_signals[0][24][12] , \s_mux2_signals[0][24][11] , 
        \s_mux2_signals[0][24][10] , \s_mux2_signals[0][24][9] , 
        \s_mux2_signals[0][24][8] , \s_mux2_signals[0][24][7] , 
        \s_mux2_signals[0][24][6] , \s_mux2_signals[0][24][5] , 
        \s_mux2_signals[0][24][4] , \s_mux2_signals[0][24][3] , 
        \s_mux2_signals[0][24][2] , \s_mux2_signals[0][24][1] , 
        \s_mux2_signals[0][24][0] }), .port1({\s_mux2_signals[0][25][31] , 
        \s_mux2_signals[0][25][30] , \s_mux2_signals[0][25][29] , 
        \s_mux2_signals[0][25][28] , \s_mux2_signals[0][25][27] , 
        \s_mux2_signals[0][25][26] , \s_mux2_signals[0][25][25] , 
        \s_mux2_signals[0][25][24] , \s_mux2_signals[0][25][23] , 
        \s_mux2_signals[0][25][22] , \s_mux2_signals[0][25][21] , 
        \s_mux2_signals[0][25][20] , \s_mux2_signals[0][25][19] , 
        \s_mux2_signals[0][25][18] , \s_mux2_signals[0][25][17] , 
        \s_mux2_signals[0][25][16] , \s_mux2_signals[0][25][15] , 
        \s_mux2_signals[0][25][14] , \s_mux2_signals[0][25][13] , 
        \s_mux2_signals[0][25][12] , \s_mux2_signals[0][25][11] , 
        \s_mux2_signals[0][25][10] , \s_mux2_signals[0][25][9] , 
        \s_mux2_signals[0][25][8] , \s_mux2_signals[0][25][7] , 
        \s_mux2_signals[0][25][6] , \s_mux2_signals[0][25][5] , 
        \s_mux2_signals[0][25][4] , \s_mux2_signals[0][25][3] , 
        \s_mux2_signals[0][25][2] , \s_mux2_signals[0][25][1] , 
        \s_mux2_signals[0][25][0] }), .sel(n26), .portY({
        \s_mux2_signals[1][24][31] , \s_mux2_signals[1][24][30] , 
        \s_mux2_signals[1][24][29] , \s_mux2_signals[1][24][28] , 
        \s_mux2_signals[1][24][27] , \s_mux2_signals[1][24][26] , 
        \s_mux2_signals[1][24][25] , \s_mux2_signals[1][24][24] , 
        \s_mux2_signals[1][24][23] , \s_mux2_signals[1][24][22] , 
        \s_mux2_signals[1][24][21] , \s_mux2_signals[1][24][20] , 
        \s_mux2_signals[1][24][19] , \s_mux2_signals[1][24][18] , 
        \s_mux2_signals[1][24][17] , \s_mux2_signals[1][24][16] , 
        \s_mux2_signals[1][24][15] , \s_mux2_signals[1][24][14] , 
        \s_mux2_signals[1][24][13] , \s_mux2_signals[1][24][12] , 
        \s_mux2_signals[1][24][11] , \s_mux2_signals[1][24][10] , 
        \s_mux2_signals[1][24][9] , \s_mux2_signals[1][24][8] , 
        \s_mux2_signals[1][24][7] , \s_mux2_signals[1][24][6] , 
        \s_mux2_signals[1][24][5] , \s_mux2_signals[1][24][4] , 
        \s_mux2_signals[1][24][3] , \s_mux2_signals[1][24][2] , 
        \s_mux2_signals[1][24][1] , \s_mux2_signals[1][24][0] }) );
  Mux_NBit_2x1_NBIT_IN32_35 MUX2_0_26 ( .port0({\s_mux2_signals[0][26][31] , 
        \s_mux2_signals[0][26][30] , \s_mux2_signals[0][26][29] , 
        \s_mux2_signals[0][26][28] , \s_mux2_signals[0][26][27] , 
        \s_mux2_signals[0][26][26] , \s_mux2_signals[0][26][25] , 
        \s_mux2_signals[0][26][24] , \s_mux2_signals[0][26][23] , 
        \s_mux2_signals[0][26][22] , \s_mux2_signals[0][26][21] , 
        \s_mux2_signals[0][26][20] , \s_mux2_signals[0][26][19] , 
        \s_mux2_signals[0][26][18] , \s_mux2_signals[0][26][17] , 
        \s_mux2_signals[0][26][16] , \s_mux2_signals[0][26][15] , 
        \s_mux2_signals[0][26][14] , \s_mux2_signals[0][26][13] , 
        \s_mux2_signals[0][26][12] , \s_mux2_signals[0][26][11] , 
        \s_mux2_signals[0][26][10] , \s_mux2_signals[0][26][9] , 
        \s_mux2_signals[0][26][8] , \s_mux2_signals[0][26][7] , 
        \s_mux2_signals[0][26][6] , \s_mux2_signals[0][26][5] , 
        \s_mux2_signals[0][26][4] , \s_mux2_signals[0][26][3] , 
        \s_mux2_signals[0][26][2] , \s_mux2_signals[0][26][1] , 
        \s_mux2_signals[0][26][0] }), .port1({\s_mux2_signals[0][27][31] , 
        \s_mux2_signals[0][27][30] , \s_mux2_signals[0][27][29] , 
        \s_mux2_signals[0][27][28] , \s_mux2_signals[0][27][27] , 
        \s_mux2_signals[0][27][26] , \s_mux2_signals[0][27][25] , 
        \s_mux2_signals[0][27][24] , \s_mux2_signals[0][27][23] , 
        \s_mux2_signals[0][27][22] , \s_mux2_signals[0][27][21] , 
        \s_mux2_signals[0][27][20] , \s_mux2_signals[0][27][19] , 
        \s_mux2_signals[0][27][18] , \s_mux2_signals[0][27][17] , 
        \s_mux2_signals[0][27][16] , \s_mux2_signals[0][27][15] , 
        \s_mux2_signals[0][27][14] , \s_mux2_signals[0][27][13] , 
        \s_mux2_signals[0][27][12] , \s_mux2_signals[0][27][11] , 
        \s_mux2_signals[0][27][10] , \s_mux2_signals[0][27][9] , 
        \s_mux2_signals[0][27][8] , \s_mux2_signals[0][27][7] , 
        \s_mux2_signals[0][27][6] , \s_mux2_signals[0][27][5] , 
        \s_mux2_signals[0][27][4] , \s_mux2_signals[0][27][3] , 
        \s_mux2_signals[0][27][2] , \s_mux2_signals[0][27][1] , 
        \s_mux2_signals[0][27][0] }), .sel(n26), .portY({
        \s_mux2_signals[1][26][31] , \s_mux2_signals[1][26][30] , 
        \s_mux2_signals[1][26][29] , \s_mux2_signals[1][26][28] , 
        \s_mux2_signals[1][26][27] , \s_mux2_signals[1][26][26] , 
        \s_mux2_signals[1][26][25] , \s_mux2_signals[1][26][24] , 
        \s_mux2_signals[1][26][23] , \s_mux2_signals[1][26][22] , 
        \s_mux2_signals[1][26][21] , \s_mux2_signals[1][26][20] , 
        \s_mux2_signals[1][26][19] , \s_mux2_signals[1][26][18] , 
        \s_mux2_signals[1][26][17] , \s_mux2_signals[1][26][16] , 
        \s_mux2_signals[1][26][15] , \s_mux2_signals[1][26][14] , 
        \s_mux2_signals[1][26][13] , \s_mux2_signals[1][26][12] , 
        \s_mux2_signals[1][26][11] , \s_mux2_signals[1][26][10] , 
        \s_mux2_signals[1][26][9] , \s_mux2_signals[1][26][8] , 
        \s_mux2_signals[1][26][7] , \s_mux2_signals[1][26][6] , 
        \s_mux2_signals[1][26][5] , \s_mux2_signals[1][26][4] , 
        \s_mux2_signals[1][26][3] , \s_mux2_signals[1][26][2] , 
        \s_mux2_signals[1][26][1] , \s_mux2_signals[1][26][0] }) );
  Mux_NBit_2x1_NBIT_IN32_34 MUX2_0_28 ( .port0({\s_mux2_signals[0][28][31] , 
        \s_mux2_signals[0][28][30] , \s_mux2_signals[0][28][29] , 
        \s_mux2_signals[0][28][28] , \s_mux2_signals[0][28][27] , 
        \s_mux2_signals[0][28][26] , \s_mux2_signals[0][28][25] , 
        \s_mux2_signals[0][28][24] , \s_mux2_signals[0][28][23] , 
        \s_mux2_signals[0][28][22] , \s_mux2_signals[0][28][21] , 
        \s_mux2_signals[0][28][20] , \s_mux2_signals[0][28][19] , 
        \s_mux2_signals[0][28][18] , \s_mux2_signals[0][28][17] , 
        \s_mux2_signals[0][28][16] , \s_mux2_signals[0][28][15] , 
        \s_mux2_signals[0][28][14] , \s_mux2_signals[0][28][13] , 
        \s_mux2_signals[0][28][12] , \s_mux2_signals[0][28][11] , 
        \s_mux2_signals[0][28][10] , \s_mux2_signals[0][28][9] , 
        \s_mux2_signals[0][28][8] , \s_mux2_signals[0][28][7] , 
        \s_mux2_signals[0][28][6] , \s_mux2_signals[0][28][5] , 
        \s_mux2_signals[0][28][4] , \s_mux2_signals[0][28][3] , 
        \s_mux2_signals[0][28][2] , \s_mux2_signals[0][28][1] , 
        \s_mux2_signals[0][28][0] }), .port1({\s_mux2_signals[0][29][31] , 
        \s_mux2_signals[0][29][30] , \s_mux2_signals[0][29][29] , 
        \s_mux2_signals[0][29][28] , \s_mux2_signals[0][29][27] , 
        \s_mux2_signals[0][29][26] , \s_mux2_signals[0][29][25] , 
        \s_mux2_signals[0][29][24] , \s_mux2_signals[0][29][23] , 
        \s_mux2_signals[0][29][22] , \s_mux2_signals[0][29][21] , 
        \s_mux2_signals[0][29][20] , \s_mux2_signals[0][29][19] , 
        \s_mux2_signals[0][29][18] , \s_mux2_signals[0][29][17] , 
        \s_mux2_signals[0][29][16] , \s_mux2_signals[0][29][15] , 
        \s_mux2_signals[0][29][14] , \s_mux2_signals[0][29][13] , 
        \s_mux2_signals[0][29][12] , \s_mux2_signals[0][29][11] , 
        \s_mux2_signals[0][29][10] , \s_mux2_signals[0][29][9] , 
        \s_mux2_signals[0][29][8] , \s_mux2_signals[0][29][7] , 
        \s_mux2_signals[0][29][6] , \s_mux2_signals[0][29][5] , 
        \s_mux2_signals[0][29][4] , \s_mux2_signals[0][29][3] , 
        \s_mux2_signals[0][29][2] , \s_mux2_signals[0][29][1] , 
        \s_mux2_signals[0][29][0] }), .sel(n27), .portY({
        \s_mux2_signals[1][28][31] , \s_mux2_signals[1][28][30] , 
        \s_mux2_signals[1][28][29] , \s_mux2_signals[1][28][28] , 
        \s_mux2_signals[1][28][27] , \s_mux2_signals[1][28][26] , 
        \s_mux2_signals[1][28][25] , \s_mux2_signals[1][28][24] , 
        \s_mux2_signals[1][28][23] , \s_mux2_signals[1][28][22] , 
        \s_mux2_signals[1][28][21] , \s_mux2_signals[1][28][20] , 
        \s_mux2_signals[1][28][19] , \s_mux2_signals[1][28][18] , 
        \s_mux2_signals[1][28][17] , \s_mux2_signals[1][28][16] , 
        \s_mux2_signals[1][28][15] , \s_mux2_signals[1][28][14] , 
        \s_mux2_signals[1][28][13] , \s_mux2_signals[1][28][12] , 
        \s_mux2_signals[1][28][11] , \s_mux2_signals[1][28][10] , 
        \s_mux2_signals[1][28][9] , \s_mux2_signals[1][28][8] , 
        \s_mux2_signals[1][28][7] , \s_mux2_signals[1][28][6] , 
        \s_mux2_signals[1][28][5] , \s_mux2_signals[1][28][4] , 
        \s_mux2_signals[1][28][3] , \s_mux2_signals[1][28][2] , 
        \s_mux2_signals[1][28][1] , \s_mux2_signals[1][28][0] }) );
  Mux_NBit_2x1_NBIT_IN32_33 MUX2_0_30 ( .port0({\s_mux2_signals[0][30][31] , 
        \s_mux2_signals[0][30][30] , \s_mux2_signals[0][30][29] , 
        \s_mux2_signals[0][30][28] , \s_mux2_signals[0][30][27] , 
        \s_mux2_signals[0][30][26] , \s_mux2_signals[0][30][25] , 
        \s_mux2_signals[0][30][24] , \s_mux2_signals[0][30][23] , 
        \s_mux2_signals[0][30][22] , \s_mux2_signals[0][30][21] , 
        \s_mux2_signals[0][30][20] , \s_mux2_signals[0][30][19] , 
        \s_mux2_signals[0][30][18] , \s_mux2_signals[0][30][17] , 
        \s_mux2_signals[0][30][16] , \s_mux2_signals[0][30][15] , 
        \s_mux2_signals[0][30][14] , \s_mux2_signals[0][30][13] , 
        \s_mux2_signals[0][30][12] , \s_mux2_signals[0][30][11] , 
        \s_mux2_signals[0][30][10] , \s_mux2_signals[0][30][9] , 
        \s_mux2_signals[0][30][8] , \s_mux2_signals[0][30][7] , 
        \s_mux2_signals[0][30][6] , \s_mux2_signals[0][30][5] , 
        \s_mux2_signals[0][30][4] , \s_mux2_signals[0][30][3] , 
        \s_mux2_signals[0][30][2] , \s_mux2_signals[0][30][1] , 
        \s_mux2_signals[0][30][0] }), .port1({\s_mux2_signals[0][31][31] , 
        \s_mux2_signals[0][31][30] , \s_mux2_signals[0][31][29] , 
        \s_mux2_signals[0][31][28] , \s_mux2_signals[0][31][27] , 
        \s_mux2_signals[0][31][26] , \s_mux2_signals[0][31][25] , 
        \s_mux2_signals[0][31][24] , \s_mux2_signals[0][31][23] , 
        \s_mux2_signals[0][31][22] , \s_mux2_signals[0][31][21] , 
        \s_mux2_signals[0][31][20] , \s_mux2_signals[0][31][19] , 
        \s_mux2_signals[0][31][18] , \s_mux2_signals[0][31][17] , 
        \s_mux2_signals[0][31][16] , \s_mux2_signals[0][31][15] , 
        \s_mux2_signals[0][31][14] , \s_mux2_signals[0][31][13] , 
        \s_mux2_signals[0][31][12] , \s_mux2_signals[0][31][11] , 
        \s_mux2_signals[0][31][10] , \s_mux2_signals[0][31][9] , 
        \s_mux2_signals[0][31][8] , \s_mux2_signals[0][31][7] , 
        \s_mux2_signals[0][31][6] , \s_mux2_signals[0][31][5] , 
        \s_mux2_signals[0][31][4] , \s_mux2_signals[0][31][3] , 
        \s_mux2_signals[0][31][2] , \s_mux2_signals[0][31][1] , n21}), .sel(
        n27), .portY({\s_mux2_signals[1][30][31] , \s_mux2_signals[1][30][30] , 
        \s_mux2_signals[1][30][29] , \s_mux2_signals[1][30][28] , 
        \s_mux2_signals[1][30][27] , \s_mux2_signals[1][30][26] , 
        \s_mux2_signals[1][30][25] , \s_mux2_signals[1][30][24] , 
        \s_mux2_signals[1][30][23] , \s_mux2_signals[1][30][22] , 
        \s_mux2_signals[1][30][21] , \s_mux2_signals[1][30][20] , 
        \s_mux2_signals[1][30][19] , \s_mux2_signals[1][30][18] , 
        \s_mux2_signals[1][30][17] , \s_mux2_signals[1][30][16] , 
        \s_mux2_signals[1][30][15] , \s_mux2_signals[1][30][14] , 
        \s_mux2_signals[1][30][13] , \s_mux2_signals[1][30][12] , 
        \s_mux2_signals[1][30][11] , \s_mux2_signals[1][30][10] , 
        \s_mux2_signals[1][30][9] , \s_mux2_signals[1][30][8] , 
        \s_mux2_signals[1][30][7] , \s_mux2_signals[1][30][6] , 
        \s_mux2_signals[1][30][5] , \s_mux2_signals[1][30][4] , 
        \s_mux2_signals[1][30][3] , \s_mux2_signals[1][30][2] , 
        \s_mux2_signals[1][30][1] , \s_mux2_signals[1][30][0] }) );
  Mux_NBit_2x1_NBIT_IN32_32 MUX2_1_0 ( .port0({\s_mux2_signals[1][0][31] , 
        \s_mux2_signals[1][0][30] , \s_mux2_signals[1][0][29] , 
        \s_mux2_signals[1][0][28] , \s_mux2_signals[1][0][27] , 
        \s_mux2_signals[1][0][26] , \s_mux2_signals[1][0][25] , 
        \s_mux2_signals[1][0][24] , \s_mux2_signals[1][0][23] , 
        \s_mux2_signals[1][0][22] , \s_mux2_signals[1][0][21] , 
        \s_mux2_signals[1][0][20] , \s_mux2_signals[1][0][19] , 
        \s_mux2_signals[1][0][18] , \s_mux2_signals[1][0][17] , 
        \s_mux2_signals[1][0][16] , \s_mux2_signals[1][0][15] , 
        \s_mux2_signals[1][0][14] , \s_mux2_signals[1][0][13] , 
        \s_mux2_signals[1][0][12] , \s_mux2_signals[1][0][11] , 
        \s_mux2_signals[1][0][10] , \s_mux2_signals[1][0][9] , 
        \s_mux2_signals[1][0][8] , \s_mux2_signals[1][0][7] , 
        \s_mux2_signals[1][0][6] , \s_mux2_signals[1][0][5] , 
        \s_mux2_signals[1][0][4] , \s_mux2_signals[1][0][3] , 
        \s_mux2_signals[1][0][2] , \s_mux2_signals[1][0][1] , 
        \s_mux2_signals[1][0][0] }), .port1({\s_mux2_signals[1][2][31] , 
        \s_mux2_signals[1][2][30] , \s_mux2_signals[1][2][29] , 
        \s_mux2_signals[1][2][28] , \s_mux2_signals[1][2][27] , 
        \s_mux2_signals[1][2][26] , \s_mux2_signals[1][2][25] , 
        \s_mux2_signals[1][2][24] , \s_mux2_signals[1][2][23] , 
        \s_mux2_signals[1][2][22] , \s_mux2_signals[1][2][21] , 
        \s_mux2_signals[1][2][20] , \s_mux2_signals[1][2][19] , 
        \s_mux2_signals[1][2][18] , \s_mux2_signals[1][2][17] , 
        \s_mux2_signals[1][2][16] , \s_mux2_signals[1][2][15] , 
        \s_mux2_signals[1][2][14] , \s_mux2_signals[1][2][13] , 
        \s_mux2_signals[1][2][12] , \s_mux2_signals[1][2][11] , 
        \s_mux2_signals[1][2][10] , \s_mux2_signals[1][2][9] , 
        \s_mux2_signals[1][2][8] , \s_mux2_signals[1][2][7] , 
        \s_mux2_signals[1][2][6] , \s_mux2_signals[1][2][5] , 
        \s_mux2_signals[1][2][4] , \s_mux2_signals[1][2][3] , 
        \s_mux2_signals[1][2][2] , \s_mux2_signals[1][2][1] , 
        \s_mux2_signals[1][2][0] }), .sel(n28), .portY({
        \s_mux2_signals[2][0][31] , \s_mux2_signals[2][0][30] , 
        \s_mux2_signals[2][0][29] , \s_mux2_signals[2][0][28] , 
        \s_mux2_signals[2][0][27] , \s_mux2_signals[2][0][26] , 
        \s_mux2_signals[2][0][25] , \s_mux2_signals[2][0][24] , 
        \s_mux2_signals[2][0][23] , \s_mux2_signals[2][0][22] , 
        \s_mux2_signals[2][0][21] , \s_mux2_signals[2][0][20] , 
        \s_mux2_signals[2][0][19] , \s_mux2_signals[2][0][18] , 
        \s_mux2_signals[2][0][17] , \s_mux2_signals[2][0][16] , 
        \s_mux2_signals[2][0][15] , \s_mux2_signals[2][0][14] , 
        \s_mux2_signals[2][0][13] , \s_mux2_signals[2][0][12] , 
        \s_mux2_signals[2][0][11] , \s_mux2_signals[2][0][10] , 
        \s_mux2_signals[2][0][9] , \s_mux2_signals[2][0][8] , 
        \s_mux2_signals[2][0][7] , \s_mux2_signals[2][0][6] , 
        \s_mux2_signals[2][0][5] , \s_mux2_signals[2][0][4] , 
        \s_mux2_signals[2][0][3] , \s_mux2_signals[2][0][2] , 
        \s_mux2_signals[2][0][1] , \s_mux2_signals[2][0][0] }) );
  Mux_NBit_2x1_NBIT_IN32_31 MUX2_1_4 ( .port0({\s_mux2_signals[1][4][31] , 
        \s_mux2_signals[1][4][30] , \s_mux2_signals[1][4][29] , 
        \s_mux2_signals[1][4][28] , \s_mux2_signals[1][4][27] , 
        \s_mux2_signals[1][4][26] , \s_mux2_signals[1][4][25] , 
        \s_mux2_signals[1][4][24] , \s_mux2_signals[1][4][23] , 
        \s_mux2_signals[1][4][22] , \s_mux2_signals[1][4][21] , 
        \s_mux2_signals[1][4][20] , \s_mux2_signals[1][4][19] , 
        \s_mux2_signals[1][4][18] , \s_mux2_signals[1][4][17] , 
        \s_mux2_signals[1][4][16] , \s_mux2_signals[1][4][15] , 
        \s_mux2_signals[1][4][14] , \s_mux2_signals[1][4][13] , 
        \s_mux2_signals[1][4][12] , \s_mux2_signals[1][4][11] , 
        \s_mux2_signals[1][4][10] , \s_mux2_signals[1][4][9] , 
        \s_mux2_signals[1][4][8] , \s_mux2_signals[1][4][7] , 
        \s_mux2_signals[1][4][6] , \s_mux2_signals[1][4][5] , 
        \s_mux2_signals[1][4][4] , \s_mux2_signals[1][4][3] , 
        \s_mux2_signals[1][4][2] , \s_mux2_signals[1][4][1] , 
        \s_mux2_signals[1][4][0] }), .port1({\s_mux2_signals[1][6][31] , 
        \s_mux2_signals[1][6][30] , \s_mux2_signals[1][6][29] , 
        \s_mux2_signals[1][6][28] , \s_mux2_signals[1][6][27] , 
        \s_mux2_signals[1][6][26] , \s_mux2_signals[1][6][25] , 
        \s_mux2_signals[1][6][24] , \s_mux2_signals[1][6][23] , 
        \s_mux2_signals[1][6][22] , \s_mux2_signals[1][6][21] , 
        \s_mux2_signals[1][6][20] , \s_mux2_signals[1][6][19] , 
        \s_mux2_signals[1][6][18] , \s_mux2_signals[1][6][17] , 
        \s_mux2_signals[1][6][16] , \s_mux2_signals[1][6][15] , 
        \s_mux2_signals[1][6][14] , \s_mux2_signals[1][6][13] , 
        \s_mux2_signals[1][6][12] , \s_mux2_signals[1][6][11] , 
        \s_mux2_signals[1][6][10] , \s_mux2_signals[1][6][9] , 
        \s_mux2_signals[1][6][8] , \s_mux2_signals[1][6][7] , 
        \s_mux2_signals[1][6][6] , \s_mux2_signals[1][6][5] , 
        \s_mux2_signals[1][6][4] , \s_mux2_signals[1][6][3] , 
        \s_mux2_signals[1][6][2] , \s_mux2_signals[1][6][1] , 
        \s_mux2_signals[1][6][0] }), .sel(n28), .portY({
        \s_mux2_signals[2][4][31] , \s_mux2_signals[2][4][30] , 
        \s_mux2_signals[2][4][29] , \s_mux2_signals[2][4][28] , 
        \s_mux2_signals[2][4][27] , \s_mux2_signals[2][4][26] , 
        \s_mux2_signals[2][4][25] , \s_mux2_signals[2][4][24] , 
        \s_mux2_signals[2][4][23] , \s_mux2_signals[2][4][22] , 
        \s_mux2_signals[2][4][21] , \s_mux2_signals[2][4][20] , 
        \s_mux2_signals[2][4][19] , \s_mux2_signals[2][4][18] , 
        \s_mux2_signals[2][4][17] , \s_mux2_signals[2][4][16] , 
        \s_mux2_signals[2][4][15] , \s_mux2_signals[2][4][14] , 
        \s_mux2_signals[2][4][13] , \s_mux2_signals[2][4][12] , 
        \s_mux2_signals[2][4][11] , \s_mux2_signals[2][4][10] , 
        \s_mux2_signals[2][4][9] , \s_mux2_signals[2][4][8] , 
        \s_mux2_signals[2][4][7] , \s_mux2_signals[2][4][6] , 
        \s_mux2_signals[2][4][5] , \s_mux2_signals[2][4][4] , 
        \s_mux2_signals[2][4][3] , \s_mux2_signals[2][4][2] , 
        \s_mux2_signals[2][4][1] , \s_mux2_signals[2][4][0] }) );
  Mux_NBit_2x1_NBIT_IN32_30 MUX2_1_8 ( .port0({\s_mux2_signals[1][8][31] , 
        \s_mux2_signals[1][8][30] , \s_mux2_signals[1][8][29] , 
        \s_mux2_signals[1][8][28] , \s_mux2_signals[1][8][27] , 
        \s_mux2_signals[1][8][26] , \s_mux2_signals[1][8][25] , 
        \s_mux2_signals[1][8][24] , \s_mux2_signals[1][8][23] , 
        \s_mux2_signals[1][8][22] , \s_mux2_signals[1][8][21] , 
        \s_mux2_signals[1][8][20] , \s_mux2_signals[1][8][19] , 
        \s_mux2_signals[1][8][18] , \s_mux2_signals[1][8][17] , 
        \s_mux2_signals[1][8][16] , \s_mux2_signals[1][8][15] , 
        \s_mux2_signals[1][8][14] , \s_mux2_signals[1][8][13] , 
        \s_mux2_signals[1][8][12] , \s_mux2_signals[1][8][11] , 
        \s_mux2_signals[1][8][10] , \s_mux2_signals[1][8][9] , 
        \s_mux2_signals[1][8][8] , \s_mux2_signals[1][8][7] , 
        \s_mux2_signals[1][8][6] , \s_mux2_signals[1][8][5] , 
        \s_mux2_signals[1][8][4] , \s_mux2_signals[1][8][3] , 
        \s_mux2_signals[1][8][2] , \s_mux2_signals[1][8][1] , 
        \s_mux2_signals[1][8][0] }), .port1({\s_mux2_signals[1][10][31] , 
        \s_mux2_signals[1][10][30] , \s_mux2_signals[1][10][29] , 
        \s_mux2_signals[1][10][28] , \s_mux2_signals[1][10][27] , 
        \s_mux2_signals[1][10][26] , \s_mux2_signals[1][10][25] , 
        \s_mux2_signals[1][10][24] , \s_mux2_signals[1][10][23] , 
        \s_mux2_signals[1][10][22] , \s_mux2_signals[1][10][21] , 
        \s_mux2_signals[1][10][20] , \s_mux2_signals[1][10][19] , 
        \s_mux2_signals[1][10][18] , \s_mux2_signals[1][10][17] , 
        \s_mux2_signals[1][10][16] , \s_mux2_signals[1][10][15] , 
        \s_mux2_signals[1][10][14] , \s_mux2_signals[1][10][13] , 
        \s_mux2_signals[1][10][12] , \s_mux2_signals[1][10][11] , 
        \s_mux2_signals[1][10][10] , \s_mux2_signals[1][10][9] , 
        \s_mux2_signals[1][10][8] , \s_mux2_signals[1][10][7] , 
        \s_mux2_signals[1][10][6] , \s_mux2_signals[1][10][5] , 
        \s_mux2_signals[1][10][4] , \s_mux2_signals[1][10][3] , 
        \s_mux2_signals[1][10][2] , \s_mux2_signals[1][10][1] , 
        \s_mux2_signals[1][10][0] }), .sel(n28), .portY({
        \s_mux2_signals[2][8][31] , \s_mux2_signals[2][8][30] , 
        \s_mux2_signals[2][8][29] , \s_mux2_signals[2][8][28] , 
        \s_mux2_signals[2][8][27] , \s_mux2_signals[2][8][26] , 
        \s_mux2_signals[2][8][25] , \s_mux2_signals[2][8][24] , 
        \s_mux2_signals[2][8][23] , \s_mux2_signals[2][8][22] , 
        \s_mux2_signals[2][8][21] , \s_mux2_signals[2][8][20] , 
        \s_mux2_signals[2][8][19] , \s_mux2_signals[2][8][18] , 
        \s_mux2_signals[2][8][17] , \s_mux2_signals[2][8][16] , 
        \s_mux2_signals[2][8][15] , \s_mux2_signals[2][8][14] , 
        \s_mux2_signals[2][8][13] , \s_mux2_signals[2][8][12] , 
        \s_mux2_signals[2][8][11] , \s_mux2_signals[2][8][10] , 
        \s_mux2_signals[2][8][9] , \s_mux2_signals[2][8][8] , 
        \s_mux2_signals[2][8][7] , \s_mux2_signals[2][8][6] , 
        \s_mux2_signals[2][8][5] , \s_mux2_signals[2][8][4] , 
        \s_mux2_signals[2][8][3] , \s_mux2_signals[2][8][2] , 
        \s_mux2_signals[2][8][1] , \s_mux2_signals[2][8][0] }) );
  Mux_NBit_2x1_NBIT_IN32_29 MUX2_1_12 ( .port0({\s_mux2_signals[1][12][31] , 
        \s_mux2_signals[1][12][30] , \s_mux2_signals[1][12][29] , 
        \s_mux2_signals[1][12][28] , \s_mux2_signals[1][12][27] , 
        \s_mux2_signals[1][12][26] , \s_mux2_signals[1][12][25] , 
        \s_mux2_signals[1][12][24] , \s_mux2_signals[1][12][23] , 
        \s_mux2_signals[1][12][22] , \s_mux2_signals[1][12][21] , 
        \s_mux2_signals[1][12][20] , \s_mux2_signals[1][12][19] , 
        \s_mux2_signals[1][12][18] , \s_mux2_signals[1][12][17] , 
        \s_mux2_signals[1][12][16] , \s_mux2_signals[1][12][15] , 
        \s_mux2_signals[1][12][14] , \s_mux2_signals[1][12][13] , 
        \s_mux2_signals[1][12][12] , \s_mux2_signals[1][12][11] , 
        \s_mux2_signals[1][12][10] , \s_mux2_signals[1][12][9] , 
        \s_mux2_signals[1][12][8] , \s_mux2_signals[1][12][7] , 
        \s_mux2_signals[1][12][6] , \s_mux2_signals[1][12][5] , 
        \s_mux2_signals[1][12][4] , \s_mux2_signals[1][12][3] , 
        \s_mux2_signals[1][12][2] , \s_mux2_signals[1][12][1] , 
        \s_mux2_signals[1][12][0] }), .port1({\s_mux2_signals[1][14][31] , 
        \s_mux2_signals[1][14][30] , \s_mux2_signals[1][14][29] , 
        \s_mux2_signals[1][14][28] , \s_mux2_signals[1][14][27] , 
        \s_mux2_signals[1][14][26] , \s_mux2_signals[1][14][25] , 
        \s_mux2_signals[1][14][24] , \s_mux2_signals[1][14][23] , 
        \s_mux2_signals[1][14][22] , \s_mux2_signals[1][14][21] , 
        \s_mux2_signals[1][14][20] , \s_mux2_signals[1][14][19] , 
        \s_mux2_signals[1][14][18] , \s_mux2_signals[1][14][17] , 
        \s_mux2_signals[1][14][16] , \s_mux2_signals[1][14][15] , 
        \s_mux2_signals[1][14][14] , \s_mux2_signals[1][14][13] , 
        \s_mux2_signals[1][14][12] , \s_mux2_signals[1][14][11] , 
        \s_mux2_signals[1][14][10] , \s_mux2_signals[1][14][9] , 
        \s_mux2_signals[1][14][8] , \s_mux2_signals[1][14][7] , 
        \s_mux2_signals[1][14][6] , \s_mux2_signals[1][14][5] , 
        \s_mux2_signals[1][14][4] , \s_mux2_signals[1][14][3] , 
        \s_mux2_signals[1][14][2] , \s_mux2_signals[1][14][1] , 
        \s_mux2_signals[1][14][0] }), .sel(n29), .portY({
        \s_mux2_signals[2][12][31] , \s_mux2_signals[2][12][30] , 
        \s_mux2_signals[2][12][29] , \s_mux2_signals[2][12][28] , 
        \s_mux2_signals[2][12][27] , \s_mux2_signals[2][12][26] , 
        \s_mux2_signals[2][12][25] , \s_mux2_signals[2][12][24] , 
        \s_mux2_signals[2][12][23] , \s_mux2_signals[2][12][22] , 
        \s_mux2_signals[2][12][21] , \s_mux2_signals[2][12][20] , 
        \s_mux2_signals[2][12][19] , \s_mux2_signals[2][12][18] , 
        \s_mux2_signals[2][12][17] , \s_mux2_signals[2][12][16] , 
        \s_mux2_signals[2][12][15] , \s_mux2_signals[2][12][14] , 
        \s_mux2_signals[2][12][13] , \s_mux2_signals[2][12][12] , 
        \s_mux2_signals[2][12][11] , \s_mux2_signals[2][12][10] , 
        \s_mux2_signals[2][12][9] , \s_mux2_signals[2][12][8] , 
        \s_mux2_signals[2][12][7] , \s_mux2_signals[2][12][6] , 
        \s_mux2_signals[2][12][5] , \s_mux2_signals[2][12][4] , 
        \s_mux2_signals[2][12][3] , \s_mux2_signals[2][12][2] , 
        \s_mux2_signals[2][12][1] , \s_mux2_signals[2][12][0] }) );
  Mux_NBit_2x1_NBIT_IN32_28 MUX2_1_16 ( .port0({\s_mux2_signals[1][16][31] , 
        \s_mux2_signals[1][16][30] , \s_mux2_signals[1][16][29] , 
        \s_mux2_signals[1][16][28] , \s_mux2_signals[1][16][27] , 
        \s_mux2_signals[1][16][26] , \s_mux2_signals[1][16][25] , 
        \s_mux2_signals[1][16][24] , \s_mux2_signals[1][16][23] , 
        \s_mux2_signals[1][16][22] , \s_mux2_signals[1][16][21] , 
        \s_mux2_signals[1][16][20] , \s_mux2_signals[1][16][19] , 
        \s_mux2_signals[1][16][18] , \s_mux2_signals[1][16][17] , 
        \s_mux2_signals[1][16][16] , \s_mux2_signals[1][16][15] , 
        \s_mux2_signals[1][16][14] , \s_mux2_signals[1][16][13] , 
        \s_mux2_signals[1][16][12] , \s_mux2_signals[1][16][11] , 
        \s_mux2_signals[1][16][10] , \s_mux2_signals[1][16][9] , 
        \s_mux2_signals[1][16][8] , \s_mux2_signals[1][16][7] , 
        \s_mux2_signals[1][16][6] , \s_mux2_signals[1][16][5] , 
        \s_mux2_signals[1][16][4] , \s_mux2_signals[1][16][3] , 
        \s_mux2_signals[1][16][2] , \s_mux2_signals[1][16][1] , 
        \s_mux2_signals[1][16][0] }), .port1({\s_mux2_signals[1][18][31] , 
        \s_mux2_signals[1][18][30] , \s_mux2_signals[1][18][29] , 
        \s_mux2_signals[1][18][28] , \s_mux2_signals[1][18][27] , 
        \s_mux2_signals[1][18][26] , \s_mux2_signals[1][18][25] , 
        \s_mux2_signals[1][18][24] , \s_mux2_signals[1][18][23] , 
        \s_mux2_signals[1][18][22] , \s_mux2_signals[1][18][21] , 
        \s_mux2_signals[1][18][20] , \s_mux2_signals[1][18][19] , 
        \s_mux2_signals[1][18][18] , \s_mux2_signals[1][18][17] , 
        \s_mux2_signals[1][18][16] , \s_mux2_signals[1][18][15] , 
        \s_mux2_signals[1][18][14] , \s_mux2_signals[1][18][13] , 
        \s_mux2_signals[1][18][12] , \s_mux2_signals[1][18][11] , 
        \s_mux2_signals[1][18][10] , \s_mux2_signals[1][18][9] , 
        \s_mux2_signals[1][18][8] , \s_mux2_signals[1][18][7] , 
        \s_mux2_signals[1][18][6] , \s_mux2_signals[1][18][5] , 
        \s_mux2_signals[1][18][4] , \s_mux2_signals[1][18][3] , 
        \s_mux2_signals[1][18][2] , \s_mux2_signals[1][18][1] , 
        \s_mux2_signals[1][18][0] }), .sel(n29), .portY({
        \s_mux2_signals[2][16][31] , \s_mux2_signals[2][16][30] , 
        \s_mux2_signals[2][16][29] , \s_mux2_signals[2][16][28] , 
        \s_mux2_signals[2][16][27] , \s_mux2_signals[2][16][26] , 
        \s_mux2_signals[2][16][25] , \s_mux2_signals[2][16][24] , 
        \s_mux2_signals[2][16][23] , \s_mux2_signals[2][16][22] , 
        \s_mux2_signals[2][16][21] , \s_mux2_signals[2][16][20] , 
        \s_mux2_signals[2][16][19] , \s_mux2_signals[2][16][18] , 
        \s_mux2_signals[2][16][17] , \s_mux2_signals[2][16][16] , 
        \s_mux2_signals[2][16][15] , \s_mux2_signals[2][16][14] , 
        \s_mux2_signals[2][16][13] , \s_mux2_signals[2][16][12] , 
        \s_mux2_signals[2][16][11] , \s_mux2_signals[2][16][10] , 
        \s_mux2_signals[2][16][9] , \s_mux2_signals[2][16][8] , 
        \s_mux2_signals[2][16][7] , \s_mux2_signals[2][16][6] , 
        \s_mux2_signals[2][16][5] , \s_mux2_signals[2][16][4] , 
        \s_mux2_signals[2][16][3] , \s_mux2_signals[2][16][2] , 
        \s_mux2_signals[2][16][1] , \s_mux2_signals[2][16][0] }) );
  Mux_NBit_2x1_NBIT_IN32_27 MUX2_1_20 ( .port0({\s_mux2_signals[1][20][31] , 
        \s_mux2_signals[1][20][30] , \s_mux2_signals[1][20][29] , 
        \s_mux2_signals[1][20][28] , \s_mux2_signals[1][20][27] , 
        \s_mux2_signals[1][20][26] , \s_mux2_signals[1][20][25] , 
        \s_mux2_signals[1][20][24] , \s_mux2_signals[1][20][23] , 
        \s_mux2_signals[1][20][22] , \s_mux2_signals[1][20][21] , 
        \s_mux2_signals[1][20][20] , \s_mux2_signals[1][20][19] , 
        \s_mux2_signals[1][20][18] , \s_mux2_signals[1][20][17] , 
        \s_mux2_signals[1][20][16] , \s_mux2_signals[1][20][15] , 
        \s_mux2_signals[1][20][14] , \s_mux2_signals[1][20][13] , 
        \s_mux2_signals[1][20][12] , \s_mux2_signals[1][20][11] , 
        \s_mux2_signals[1][20][10] , \s_mux2_signals[1][20][9] , 
        \s_mux2_signals[1][20][8] , \s_mux2_signals[1][20][7] , 
        \s_mux2_signals[1][20][6] , \s_mux2_signals[1][20][5] , 
        \s_mux2_signals[1][20][4] , \s_mux2_signals[1][20][3] , 
        \s_mux2_signals[1][20][2] , \s_mux2_signals[1][20][1] , 
        \s_mux2_signals[1][20][0] }), .port1({\s_mux2_signals[1][22][31] , 
        \s_mux2_signals[1][22][30] , \s_mux2_signals[1][22][29] , 
        \s_mux2_signals[1][22][28] , \s_mux2_signals[1][22][27] , 
        \s_mux2_signals[1][22][26] , \s_mux2_signals[1][22][25] , 
        \s_mux2_signals[1][22][24] , \s_mux2_signals[1][22][23] , 
        \s_mux2_signals[1][22][22] , \s_mux2_signals[1][22][21] , 
        \s_mux2_signals[1][22][20] , \s_mux2_signals[1][22][19] , 
        \s_mux2_signals[1][22][18] , \s_mux2_signals[1][22][17] , 
        \s_mux2_signals[1][22][16] , \s_mux2_signals[1][22][15] , 
        \s_mux2_signals[1][22][14] , \s_mux2_signals[1][22][13] , 
        \s_mux2_signals[1][22][12] , \s_mux2_signals[1][22][11] , 
        \s_mux2_signals[1][22][10] , \s_mux2_signals[1][22][9] , 
        \s_mux2_signals[1][22][8] , \s_mux2_signals[1][22][7] , 
        \s_mux2_signals[1][22][6] , \s_mux2_signals[1][22][5] , 
        \s_mux2_signals[1][22][4] , \s_mux2_signals[1][22][3] , 
        \s_mux2_signals[1][22][2] , \s_mux2_signals[1][22][1] , 
        \s_mux2_signals[1][22][0] }), .sel(n29), .portY({
        \s_mux2_signals[2][20][31] , \s_mux2_signals[2][20][30] , 
        \s_mux2_signals[2][20][29] , \s_mux2_signals[2][20][28] , 
        \s_mux2_signals[2][20][27] , \s_mux2_signals[2][20][26] , 
        \s_mux2_signals[2][20][25] , \s_mux2_signals[2][20][24] , 
        \s_mux2_signals[2][20][23] , \s_mux2_signals[2][20][22] , 
        \s_mux2_signals[2][20][21] , \s_mux2_signals[2][20][20] , 
        \s_mux2_signals[2][20][19] , \s_mux2_signals[2][20][18] , 
        \s_mux2_signals[2][20][17] , \s_mux2_signals[2][20][16] , 
        \s_mux2_signals[2][20][15] , \s_mux2_signals[2][20][14] , 
        \s_mux2_signals[2][20][13] , \s_mux2_signals[2][20][12] , 
        \s_mux2_signals[2][20][11] , \s_mux2_signals[2][20][10] , 
        \s_mux2_signals[2][20][9] , \s_mux2_signals[2][20][8] , 
        \s_mux2_signals[2][20][7] , \s_mux2_signals[2][20][6] , 
        \s_mux2_signals[2][20][5] , \s_mux2_signals[2][20][4] , 
        \s_mux2_signals[2][20][3] , \s_mux2_signals[2][20][2] , 
        \s_mux2_signals[2][20][1] , \s_mux2_signals[2][20][0] }) );
  Mux_NBit_2x1_NBIT_IN32_26 MUX2_1_24 ( .port0({\s_mux2_signals[1][24][31] , 
        \s_mux2_signals[1][24][30] , \s_mux2_signals[1][24][29] , 
        \s_mux2_signals[1][24][28] , \s_mux2_signals[1][24][27] , 
        \s_mux2_signals[1][24][26] , \s_mux2_signals[1][24][25] , 
        \s_mux2_signals[1][24][24] , \s_mux2_signals[1][24][23] , 
        \s_mux2_signals[1][24][22] , \s_mux2_signals[1][24][21] , 
        \s_mux2_signals[1][24][20] , \s_mux2_signals[1][24][19] , 
        \s_mux2_signals[1][24][18] , \s_mux2_signals[1][24][17] , 
        \s_mux2_signals[1][24][16] , \s_mux2_signals[1][24][15] , 
        \s_mux2_signals[1][24][14] , \s_mux2_signals[1][24][13] , 
        \s_mux2_signals[1][24][12] , \s_mux2_signals[1][24][11] , 
        \s_mux2_signals[1][24][10] , \s_mux2_signals[1][24][9] , 
        \s_mux2_signals[1][24][8] , \s_mux2_signals[1][24][7] , 
        \s_mux2_signals[1][24][6] , \s_mux2_signals[1][24][5] , 
        \s_mux2_signals[1][24][4] , \s_mux2_signals[1][24][3] , 
        \s_mux2_signals[1][24][2] , \s_mux2_signals[1][24][1] , 
        \s_mux2_signals[1][24][0] }), .port1({\s_mux2_signals[1][26][31] , 
        \s_mux2_signals[1][26][30] , \s_mux2_signals[1][26][29] , 
        \s_mux2_signals[1][26][28] , \s_mux2_signals[1][26][27] , 
        \s_mux2_signals[1][26][26] , \s_mux2_signals[1][26][25] , 
        \s_mux2_signals[1][26][24] , \s_mux2_signals[1][26][23] , 
        \s_mux2_signals[1][26][22] , \s_mux2_signals[1][26][21] , 
        \s_mux2_signals[1][26][20] , \s_mux2_signals[1][26][19] , 
        \s_mux2_signals[1][26][18] , \s_mux2_signals[1][26][17] , 
        \s_mux2_signals[1][26][16] , \s_mux2_signals[1][26][15] , 
        \s_mux2_signals[1][26][14] , \s_mux2_signals[1][26][13] , 
        \s_mux2_signals[1][26][12] , \s_mux2_signals[1][26][11] , 
        \s_mux2_signals[1][26][10] , \s_mux2_signals[1][26][9] , 
        \s_mux2_signals[1][26][8] , \s_mux2_signals[1][26][7] , 
        \s_mux2_signals[1][26][6] , \s_mux2_signals[1][26][5] , 
        \s_mux2_signals[1][26][4] , \s_mux2_signals[1][26][3] , 
        \s_mux2_signals[1][26][2] , \s_mux2_signals[1][26][1] , 
        \s_mux2_signals[1][26][0] }), .sel(n30), .portY({
        \s_mux2_signals[2][24][31] , \s_mux2_signals[2][24][30] , 
        \s_mux2_signals[2][24][29] , \s_mux2_signals[2][24][28] , 
        \s_mux2_signals[2][24][27] , \s_mux2_signals[2][24][26] , 
        \s_mux2_signals[2][24][25] , \s_mux2_signals[2][24][24] , 
        \s_mux2_signals[2][24][23] , \s_mux2_signals[2][24][22] , 
        \s_mux2_signals[2][24][21] , \s_mux2_signals[2][24][20] , 
        \s_mux2_signals[2][24][19] , \s_mux2_signals[2][24][18] , 
        \s_mux2_signals[2][24][17] , \s_mux2_signals[2][24][16] , 
        \s_mux2_signals[2][24][15] , \s_mux2_signals[2][24][14] , 
        \s_mux2_signals[2][24][13] , \s_mux2_signals[2][24][12] , 
        \s_mux2_signals[2][24][11] , \s_mux2_signals[2][24][10] , 
        \s_mux2_signals[2][24][9] , \s_mux2_signals[2][24][8] , 
        \s_mux2_signals[2][24][7] , \s_mux2_signals[2][24][6] , 
        \s_mux2_signals[2][24][5] , \s_mux2_signals[2][24][4] , 
        \s_mux2_signals[2][24][3] , \s_mux2_signals[2][24][2] , 
        \s_mux2_signals[2][24][1] , \s_mux2_signals[2][24][0] }) );
  Mux_NBit_2x1_NBIT_IN32_25 MUX2_1_28 ( .port0({\s_mux2_signals[1][28][31] , 
        \s_mux2_signals[1][28][30] , \s_mux2_signals[1][28][29] , 
        \s_mux2_signals[1][28][28] , \s_mux2_signals[1][28][27] , 
        \s_mux2_signals[1][28][26] , \s_mux2_signals[1][28][25] , 
        \s_mux2_signals[1][28][24] , \s_mux2_signals[1][28][23] , 
        \s_mux2_signals[1][28][22] , \s_mux2_signals[1][28][21] , 
        \s_mux2_signals[1][28][20] , \s_mux2_signals[1][28][19] , 
        \s_mux2_signals[1][28][18] , \s_mux2_signals[1][28][17] , 
        \s_mux2_signals[1][28][16] , \s_mux2_signals[1][28][15] , 
        \s_mux2_signals[1][28][14] , \s_mux2_signals[1][28][13] , 
        \s_mux2_signals[1][28][12] , \s_mux2_signals[1][28][11] , 
        \s_mux2_signals[1][28][10] , \s_mux2_signals[1][28][9] , 
        \s_mux2_signals[1][28][8] , \s_mux2_signals[1][28][7] , 
        \s_mux2_signals[1][28][6] , \s_mux2_signals[1][28][5] , 
        \s_mux2_signals[1][28][4] , \s_mux2_signals[1][28][3] , 
        \s_mux2_signals[1][28][2] , \s_mux2_signals[1][28][1] , 
        \s_mux2_signals[1][28][0] }), .port1({\s_mux2_signals[1][30][31] , 
        \s_mux2_signals[1][30][30] , \s_mux2_signals[1][30][29] , 
        \s_mux2_signals[1][30][28] , \s_mux2_signals[1][30][27] , 
        \s_mux2_signals[1][30][26] , \s_mux2_signals[1][30][25] , 
        \s_mux2_signals[1][30][24] , \s_mux2_signals[1][30][23] , 
        \s_mux2_signals[1][30][22] , \s_mux2_signals[1][30][21] , 
        \s_mux2_signals[1][30][20] , \s_mux2_signals[1][30][19] , 
        \s_mux2_signals[1][30][18] , \s_mux2_signals[1][30][17] , 
        \s_mux2_signals[1][30][16] , \s_mux2_signals[1][30][15] , 
        \s_mux2_signals[1][30][14] , \s_mux2_signals[1][30][13] , 
        \s_mux2_signals[1][30][12] , \s_mux2_signals[1][30][11] , 
        \s_mux2_signals[1][30][10] , \s_mux2_signals[1][30][9] , 
        \s_mux2_signals[1][30][8] , \s_mux2_signals[1][30][7] , 
        \s_mux2_signals[1][30][6] , \s_mux2_signals[1][30][5] , 
        \s_mux2_signals[1][30][4] , \s_mux2_signals[1][30][3] , 
        \s_mux2_signals[1][30][2] , \s_mux2_signals[1][30][1] , 
        \s_mux2_signals[1][30][0] }), .sel(n30), .portY({
        \s_mux2_signals[2][28][31] , \s_mux2_signals[2][28][30] , 
        \s_mux2_signals[2][28][29] , \s_mux2_signals[2][28][28] , 
        \s_mux2_signals[2][28][27] , \s_mux2_signals[2][28][26] , 
        \s_mux2_signals[2][28][25] , \s_mux2_signals[2][28][24] , 
        \s_mux2_signals[2][28][23] , \s_mux2_signals[2][28][22] , 
        \s_mux2_signals[2][28][21] , \s_mux2_signals[2][28][20] , 
        \s_mux2_signals[2][28][19] , \s_mux2_signals[2][28][18] , 
        \s_mux2_signals[2][28][17] , \s_mux2_signals[2][28][16] , 
        \s_mux2_signals[2][28][15] , \s_mux2_signals[2][28][14] , 
        \s_mux2_signals[2][28][13] , \s_mux2_signals[2][28][12] , 
        \s_mux2_signals[2][28][11] , \s_mux2_signals[2][28][10] , 
        \s_mux2_signals[2][28][9] , \s_mux2_signals[2][28][8] , 
        \s_mux2_signals[2][28][7] , \s_mux2_signals[2][28][6] , 
        \s_mux2_signals[2][28][5] , \s_mux2_signals[2][28][4] , 
        \s_mux2_signals[2][28][3] , \s_mux2_signals[2][28][2] , 
        \s_mux2_signals[2][28][1] , \s_mux2_signals[2][28][0] }) );
  Mux_NBit_2x1_NBIT_IN32_24 MUX2_2_0 ( .port0({\s_mux2_signals[2][0][31] , 
        \s_mux2_signals[2][0][30] , \s_mux2_signals[2][0][29] , 
        \s_mux2_signals[2][0][28] , \s_mux2_signals[2][0][27] , 
        \s_mux2_signals[2][0][26] , \s_mux2_signals[2][0][25] , 
        \s_mux2_signals[2][0][24] , \s_mux2_signals[2][0][23] , 
        \s_mux2_signals[2][0][22] , \s_mux2_signals[2][0][21] , 
        \s_mux2_signals[2][0][20] , \s_mux2_signals[2][0][19] , 
        \s_mux2_signals[2][0][18] , \s_mux2_signals[2][0][17] , 
        \s_mux2_signals[2][0][16] , \s_mux2_signals[2][0][15] , 
        \s_mux2_signals[2][0][14] , \s_mux2_signals[2][0][13] , 
        \s_mux2_signals[2][0][12] , \s_mux2_signals[2][0][11] , 
        \s_mux2_signals[2][0][10] , \s_mux2_signals[2][0][9] , 
        \s_mux2_signals[2][0][8] , \s_mux2_signals[2][0][7] , 
        \s_mux2_signals[2][0][6] , \s_mux2_signals[2][0][5] , 
        \s_mux2_signals[2][0][4] , \s_mux2_signals[2][0][3] , 
        \s_mux2_signals[2][0][2] , \s_mux2_signals[2][0][1] , 
        \s_mux2_signals[2][0][0] }), .port1({\s_mux2_signals[2][4][31] , 
        \s_mux2_signals[2][4][30] , \s_mux2_signals[2][4][29] , 
        \s_mux2_signals[2][4][28] , \s_mux2_signals[2][4][27] , 
        \s_mux2_signals[2][4][26] , \s_mux2_signals[2][4][25] , 
        \s_mux2_signals[2][4][24] , \s_mux2_signals[2][4][23] , 
        \s_mux2_signals[2][4][22] , \s_mux2_signals[2][4][21] , 
        \s_mux2_signals[2][4][20] , \s_mux2_signals[2][4][19] , 
        \s_mux2_signals[2][4][18] , \s_mux2_signals[2][4][17] , 
        \s_mux2_signals[2][4][16] , \s_mux2_signals[2][4][15] , 
        \s_mux2_signals[2][4][14] , \s_mux2_signals[2][4][13] , 
        \s_mux2_signals[2][4][12] , \s_mux2_signals[2][4][11] , 
        \s_mux2_signals[2][4][10] , \s_mux2_signals[2][4][9] , 
        \s_mux2_signals[2][4][8] , \s_mux2_signals[2][4][7] , 
        \s_mux2_signals[2][4][6] , \s_mux2_signals[2][4][5] , 
        \s_mux2_signals[2][4][4] , \s_mux2_signals[2][4][3] , 
        \s_mux2_signals[2][4][2] , \s_mux2_signals[2][4][1] , 
        \s_mux2_signals[2][4][0] }), .sel(n31), .portY({
        \s_mux2_signals[3][0][31] , \s_mux2_signals[3][0][30] , 
        \s_mux2_signals[3][0][29] , \s_mux2_signals[3][0][28] , 
        \s_mux2_signals[3][0][27] , \s_mux2_signals[3][0][26] , 
        \s_mux2_signals[3][0][25] , \s_mux2_signals[3][0][24] , 
        \s_mux2_signals[3][0][23] , \s_mux2_signals[3][0][22] , 
        \s_mux2_signals[3][0][21] , \s_mux2_signals[3][0][20] , 
        \s_mux2_signals[3][0][19] , \s_mux2_signals[3][0][18] , 
        \s_mux2_signals[3][0][17] , \s_mux2_signals[3][0][16] , 
        \s_mux2_signals[3][0][15] , \s_mux2_signals[3][0][14] , 
        \s_mux2_signals[3][0][13] , \s_mux2_signals[3][0][12] , 
        \s_mux2_signals[3][0][11] , \s_mux2_signals[3][0][10] , 
        \s_mux2_signals[3][0][9] , \s_mux2_signals[3][0][8] , 
        \s_mux2_signals[3][0][7] , \s_mux2_signals[3][0][6] , 
        \s_mux2_signals[3][0][5] , \s_mux2_signals[3][0][4] , 
        \s_mux2_signals[3][0][3] , \s_mux2_signals[3][0][2] , 
        \s_mux2_signals[3][0][1] , \s_mux2_signals[3][0][0] }) );
  Mux_NBit_2x1_NBIT_IN32_23 MUX2_2_8 ( .port0({\s_mux2_signals[2][8][31] , 
        \s_mux2_signals[2][8][30] , \s_mux2_signals[2][8][29] , 
        \s_mux2_signals[2][8][28] , \s_mux2_signals[2][8][27] , 
        \s_mux2_signals[2][8][26] , \s_mux2_signals[2][8][25] , 
        \s_mux2_signals[2][8][24] , \s_mux2_signals[2][8][23] , 
        \s_mux2_signals[2][8][22] , \s_mux2_signals[2][8][21] , 
        \s_mux2_signals[2][8][20] , \s_mux2_signals[2][8][19] , 
        \s_mux2_signals[2][8][18] , \s_mux2_signals[2][8][17] , 
        \s_mux2_signals[2][8][16] , \s_mux2_signals[2][8][15] , 
        \s_mux2_signals[2][8][14] , \s_mux2_signals[2][8][13] , 
        \s_mux2_signals[2][8][12] , \s_mux2_signals[2][8][11] , 
        \s_mux2_signals[2][8][10] , \s_mux2_signals[2][8][9] , 
        \s_mux2_signals[2][8][8] , \s_mux2_signals[2][8][7] , 
        \s_mux2_signals[2][8][6] , \s_mux2_signals[2][8][5] , 
        \s_mux2_signals[2][8][4] , \s_mux2_signals[2][8][3] , 
        \s_mux2_signals[2][8][2] , \s_mux2_signals[2][8][1] , 
        \s_mux2_signals[2][8][0] }), .port1({\s_mux2_signals[2][12][31] , 
        \s_mux2_signals[2][12][30] , \s_mux2_signals[2][12][29] , 
        \s_mux2_signals[2][12][28] , \s_mux2_signals[2][12][27] , 
        \s_mux2_signals[2][12][26] , \s_mux2_signals[2][12][25] , 
        \s_mux2_signals[2][12][24] , \s_mux2_signals[2][12][23] , 
        \s_mux2_signals[2][12][22] , \s_mux2_signals[2][12][21] , 
        \s_mux2_signals[2][12][20] , \s_mux2_signals[2][12][19] , 
        \s_mux2_signals[2][12][18] , \s_mux2_signals[2][12][17] , 
        \s_mux2_signals[2][12][16] , \s_mux2_signals[2][12][15] , 
        \s_mux2_signals[2][12][14] , \s_mux2_signals[2][12][13] , 
        \s_mux2_signals[2][12][12] , \s_mux2_signals[2][12][11] , 
        \s_mux2_signals[2][12][10] , \s_mux2_signals[2][12][9] , 
        \s_mux2_signals[2][12][8] , \s_mux2_signals[2][12][7] , 
        \s_mux2_signals[2][12][6] , \s_mux2_signals[2][12][5] , 
        \s_mux2_signals[2][12][4] , \s_mux2_signals[2][12][3] , 
        \s_mux2_signals[2][12][2] , \s_mux2_signals[2][12][1] , 
        \s_mux2_signals[2][12][0] }), .sel(n31), .portY({
        \s_mux2_signals[3][8][31] , \s_mux2_signals[3][8][30] , 
        \s_mux2_signals[3][8][29] , \s_mux2_signals[3][8][28] , 
        \s_mux2_signals[3][8][27] , \s_mux2_signals[3][8][26] , 
        \s_mux2_signals[3][8][25] , \s_mux2_signals[3][8][24] , 
        \s_mux2_signals[3][8][23] , \s_mux2_signals[3][8][22] , 
        \s_mux2_signals[3][8][21] , \s_mux2_signals[3][8][20] , 
        \s_mux2_signals[3][8][19] , \s_mux2_signals[3][8][18] , 
        \s_mux2_signals[3][8][17] , \s_mux2_signals[3][8][16] , 
        \s_mux2_signals[3][8][15] , \s_mux2_signals[3][8][14] , 
        \s_mux2_signals[3][8][13] , \s_mux2_signals[3][8][12] , 
        \s_mux2_signals[3][8][11] , \s_mux2_signals[3][8][10] , 
        \s_mux2_signals[3][8][9] , \s_mux2_signals[3][8][8] , 
        \s_mux2_signals[3][8][7] , \s_mux2_signals[3][8][6] , 
        \s_mux2_signals[3][8][5] , \s_mux2_signals[3][8][4] , 
        \s_mux2_signals[3][8][3] , \s_mux2_signals[3][8][2] , 
        \s_mux2_signals[3][8][1] , \s_mux2_signals[3][8][0] }) );
  Mux_NBit_2x1_NBIT_IN32_22 MUX2_2_16 ( .port0({\s_mux2_signals[2][16][31] , 
        \s_mux2_signals[2][16][30] , \s_mux2_signals[2][16][29] , 
        \s_mux2_signals[2][16][28] , \s_mux2_signals[2][16][27] , 
        \s_mux2_signals[2][16][26] , \s_mux2_signals[2][16][25] , 
        \s_mux2_signals[2][16][24] , \s_mux2_signals[2][16][23] , 
        \s_mux2_signals[2][16][22] , \s_mux2_signals[2][16][21] , 
        \s_mux2_signals[2][16][20] , \s_mux2_signals[2][16][19] , 
        \s_mux2_signals[2][16][18] , \s_mux2_signals[2][16][17] , 
        \s_mux2_signals[2][16][16] , \s_mux2_signals[2][16][15] , 
        \s_mux2_signals[2][16][14] , \s_mux2_signals[2][16][13] , 
        \s_mux2_signals[2][16][12] , \s_mux2_signals[2][16][11] , 
        \s_mux2_signals[2][16][10] , \s_mux2_signals[2][16][9] , 
        \s_mux2_signals[2][16][8] , \s_mux2_signals[2][16][7] , 
        \s_mux2_signals[2][16][6] , \s_mux2_signals[2][16][5] , 
        \s_mux2_signals[2][16][4] , \s_mux2_signals[2][16][3] , 
        \s_mux2_signals[2][16][2] , \s_mux2_signals[2][16][1] , 
        \s_mux2_signals[2][16][0] }), .port1({\s_mux2_signals[2][20][31] , 
        \s_mux2_signals[2][20][30] , \s_mux2_signals[2][20][29] , 
        \s_mux2_signals[2][20][28] , \s_mux2_signals[2][20][27] , 
        \s_mux2_signals[2][20][26] , \s_mux2_signals[2][20][25] , 
        \s_mux2_signals[2][20][24] , \s_mux2_signals[2][20][23] , 
        \s_mux2_signals[2][20][22] , \s_mux2_signals[2][20][21] , 
        \s_mux2_signals[2][20][20] , \s_mux2_signals[2][20][19] , 
        \s_mux2_signals[2][20][18] , \s_mux2_signals[2][20][17] , 
        \s_mux2_signals[2][20][16] , \s_mux2_signals[2][20][15] , 
        \s_mux2_signals[2][20][14] , \s_mux2_signals[2][20][13] , 
        \s_mux2_signals[2][20][12] , \s_mux2_signals[2][20][11] , 
        \s_mux2_signals[2][20][10] , \s_mux2_signals[2][20][9] , 
        \s_mux2_signals[2][20][8] , \s_mux2_signals[2][20][7] , 
        \s_mux2_signals[2][20][6] , \s_mux2_signals[2][20][5] , 
        \s_mux2_signals[2][20][4] , \s_mux2_signals[2][20][3] , 
        \s_mux2_signals[2][20][2] , \s_mux2_signals[2][20][1] , 
        \s_mux2_signals[2][20][0] }), .sel(n31), .portY({
        \s_mux2_signals[3][16][31] , \s_mux2_signals[3][16][30] , 
        \s_mux2_signals[3][16][29] , \s_mux2_signals[3][16][28] , 
        \s_mux2_signals[3][16][27] , \s_mux2_signals[3][16][26] , 
        \s_mux2_signals[3][16][25] , \s_mux2_signals[3][16][24] , 
        \s_mux2_signals[3][16][23] , \s_mux2_signals[3][16][22] , 
        \s_mux2_signals[3][16][21] , \s_mux2_signals[3][16][20] , 
        \s_mux2_signals[3][16][19] , \s_mux2_signals[3][16][18] , 
        \s_mux2_signals[3][16][17] , \s_mux2_signals[3][16][16] , 
        \s_mux2_signals[3][16][15] , \s_mux2_signals[3][16][14] , 
        \s_mux2_signals[3][16][13] , \s_mux2_signals[3][16][12] , 
        \s_mux2_signals[3][16][11] , \s_mux2_signals[3][16][10] , 
        \s_mux2_signals[3][16][9] , \s_mux2_signals[3][16][8] , 
        \s_mux2_signals[3][16][7] , \s_mux2_signals[3][16][6] , 
        \s_mux2_signals[3][16][5] , \s_mux2_signals[3][16][4] , 
        \s_mux2_signals[3][16][3] , \s_mux2_signals[3][16][2] , 
        \s_mux2_signals[3][16][1] , \s_mux2_signals[3][16][0] }) );
  Mux_NBit_2x1_NBIT_IN32_21 MUX2_2_24 ( .port0({\s_mux2_signals[2][24][31] , 
        \s_mux2_signals[2][24][30] , \s_mux2_signals[2][24][29] , 
        \s_mux2_signals[2][24][28] , \s_mux2_signals[2][24][27] , 
        \s_mux2_signals[2][24][26] , \s_mux2_signals[2][24][25] , 
        \s_mux2_signals[2][24][24] , \s_mux2_signals[2][24][23] , 
        \s_mux2_signals[2][24][22] , \s_mux2_signals[2][24][21] , 
        \s_mux2_signals[2][24][20] , \s_mux2_signals[2][24][19] , 
        \s_mux2_signals[2][24][18] , \s_mux2_signals[2][24][17] , 
        \s_mux2_signals[2][24][16] , \s_mux2_signals[2][24][15] , 
        \s_mux2_signals[2][24][14] , \s_mux2_signals[2][24][13] , 
        \s_mux2_signals[2][24][12] , \s_mux2_signals[2][24][11] , 
        \s_mux2_signals[2][24][10] , \s_mux2_signals[2][24][9] , 
        \s_mux2_signals[2][24][8] , \s_mux2_signals[2][24][7] , 
        \s_mux2_signals[2][24][6] , \s_mux2_signals[2][24][5] , 
        \s_mux2_signals[2][24][4] , \s_mux2_signals[2][24][3] , 
        \s_mux2_signals[2][24][2] , \s_mux2_signals[2][24][1] , 
        \s_mux2_signals[2][24][0] }), .port1({\s_mux2_signals[2][28][31] , 
        \s_mux2_signals[2][28][30] , \s_mux2_signals[2][28][29] , 
        \s_mux2_signals[2][28][28] , \s_mux2_signals[2][28][27] , 
        \s_mux2_signals[2][28][26] , \s_mux2_signals[2][28][25] , 
        \s_mux2_signals[2][28][24] , \s_mux2_signals[2][28][23] , 
        \s_mux2_signals[2][28][22] , \s_mux2_signals[2][28][21] , 
        \s_mux2_signals[2][28][20] , \s_mux2_signals[2][28][19] , 
        \s_mux2_signals[2][28][18] , \s_mux2_signals[2][28][17] , 
        \s_mux2_signals[2][28][16] , \s_mux2_signals[2][28][15] , 
        \s_mux2_signals[2][28][14] , \s_mux2_signals[2][28][13] , 
        \s_mux2_signals[2][28][12] , \s_mux2_signals[2][28][11] , 
        \s_mux2_signals[2][28][10] , \s_mux2_signals[2][28][9] , 
        \s_mux2_signals[2][28][8] , \s_mux2_signals[2][28][7] , 
        \s_mux2_signals[2][28][6] , \s_mux2_signals[2][28][5] , 
        \s_mux2_signals[2][28][4] , \s_mux2_signals[2][28][3] , 
        \s_mux2_signals[2][28][2] , \s_mux2_signals[2][28][1] , 
        \s_mux2_signals[2][28][0] }), .sel(n31), .portY({
        \s_mux2_signals[3][24][31] , \s_mux2_signals[3][24][30] , 
        \s_mux2_signals[3][24][29] , \s_mux2_signals[3][24][28] , 
        \s_mux2_signals[3][24][27] , \s_mux2_signals[3][24][26] , 
        \s_mux2_signals[3][24][25] , \s_mux2_signals[3][24][24] , 
        \s_mux2_signals[3][24][23] , \s_mux2_signals[3][24][22] , 
        \s_mux2_signals[3][24][21] , \s_mux2_signals[3][24][20] , 
        \s_mux2_signals[3][24][19] , \s_mux2_signals[3][24][18] , 
        \s_mux2_signals[3][24][17] , \s_mux2_signals[3][24][16] , 
        \s_mux2_signals[3][24][15] , \s_mux2_signals[3][24][14] , 
        \s_mux2_signals[3][24][13] , \s_mux2_signals[3][24][12] , 
        \s_mux2_signals[3][24][11] , \s_mux2_signals[3][24][10] , 
        \s_mux2_signals[3][24][9] , \s_mux2_signals[3][24][8] , 
        \s_mux2_signals[3][24][7] , \s_mux2_signals[3][24][6] , 
        \s_mux2_signals[3][24][5] , \s_mux2_signals[3][24][4] , 
        \s_mux2_signals[3][24][3] , \s_mux2_signals[3][24][2] , 
        \s_mux2_signals[3][24][1] , \s_mux2_signals[3][24][0] }) );
  Mux_NBit_2x1_NBIT_IN32_20 MUX2_3_0 ( .port0({\s_mux2_signals[3][0][31] , 
        \s_mux2_signals[3][0][30] , \s_mux2_signals[3][0][29] , 
        \s_mux2_signals[3][0][28] , \s_mux2_signals[3][0][27] , 
        \s_mux2_signals[3][0][26] , \s_mux2_signals[3][0][25] , 
        \s_mux2_signals[3][0][24] , \s_mux2_signals[3][0][23] , 
        \s_mux2_signals[3][0][22] , \s_mux2_signals[3][0][21] , 
        \s_mux2_signals[3][0][20] , \s_mux2_signals[3][0][19] , 
        \s_mux2_signals[3][0][18] , \s_mux2_signals[3][0][17] , 
        \s_mux2_signals[3][0][16] , \s_mux2_signals[3][0][15] , 
        \s_mux2_signals[3][0][14] , \s_mux2_signals[3][0][13] , 
        \s_mux2_signals[3][0][12] , \s_mux2_signals[3][0][11] , 
        \s_mux2_signals[3][0][10] , \s_mux2_signals[3][0][9] , 
        \s_mux2_signals[3][0][8] , \s_mux2_signals[3][0][7] , 
        \s_mux2_signals[3][0][6] , \s_mux2_signals[3][0][5] , 
        \s_mux2_signals[3][0][4] , \s_mux2_signals[3][0][3] , 
        \s_mux2_signals[3][0][2] , \s_mux2_signals[3][0][1] , 
        \s_mux2_signals[3][0][0] }), .port1({\s_mux2_signals[3][8][31] , 
        \s_mux2_signals[3][8][30] , \s_mux2_signals[3][8][29] , 
        \s_mux2_signals[3][8][28] , \s_mux2_signals[3][8][27] , 
        \s_mux2_signals[3][8][26] , \s_mux2_signals[3][8][25] , 
        \s_mux2_signals[3][8][24] , \s_mux2_signals[3][8][23] , 
        \s_mux2_signals[3][8][22] , \s_mux2_signals[3][8][21] , 
        \s_mux2_signals[3][8][20] , \s_mux2_signals[3][8][19] , 
        \s_mux2_signals[3][8][18] , \s_mux2_signals[3][8][17] , 
        \s_mux2_signals[3][8][16] , \s_mux2_signals[3][8][15] , 
        \s_mux2_signals[3][8][14] , \s_mux2_signals[3][8][13] , 
        \s_mux2_signals[3][8][12] , \s_mux2_signals[3][8][11] , 
        \s_mux2_signals[3][8][10] , \s_mux2_signals[3][8][9] , 
        \s_mux2_signals[3][8][8] , \s_mux2_signals[3][8][7] , 
        \s_mux2_signals[3][8][6] , \s_mux2_signals[3][8][5] , 
        \s_mux2_signals[3][8][4] , \s_mux2_signals[3][8][3] , 
        \s_mux2_signals[3][8][2] , \s_mux2_signals[3][8][1] , 
        \s_mux2_signals[3][8][0] }), .sel(s_addrRd2_Fei_Tmux[3]), .portY({
        \s_mux2_signals[4][0][31] , \s_mux2_signals[4][0][30] , 
        \s_mux2_signals[4][0][29] , \s_mux2_signals[4][0][28] , 
        \s_mux2_signals[4][0][27] , \s_mux2_signals[4][0][26] , 
        \s_mux2_signals[4][0][25] , \s_mux2_signals[4][0][24] , 
        \s_mux2_signals[4][0][23] , \s_mux2_signals[4][0][22] , 
        \s_mux2_signals[4][0][21] , \s_mux2_signals[4][0][20] , 
        \s_mux2_signals[4][0][19] , \s_mux2_signals[4][0][18] , 
        \s_mux2_signals[4][0][17] , \s_mux2_signals[4][0][16] , 
        \s_mux2_signals[4][0][15] , \s_mux2_signals[4][0][14] , 
        \s_mux2_signals[4][0][13] , \s_mux2_signals[4][0][12] , 
        \s_mux2_signals[4][0][11] , \s_mux2_signals[4][0][10] , 
        \s_mux2_signals[4][0][9] , \s_mux2_signals[4][0][8] , 
        \s_mux2_signals[4][0][7] , \s_mux2_signals[4][0][6] , 
        \s_mux2_signals[4][0][5] , \s_mux2_signals[4][0][4] , 
        \s_mux2_signals[4][0][3] , \s_mux2_signals[4][0][2] , 
        \s_mux2_signals[4][0][1] , \s_mux2_signals[4][0][0] }) );
  Mux_NBit_2x1_NBIT_IN32_19 MUX2_3_16 ( .port0({\s_mux2_signals[3][16][31] , 
        \s_mux2_signals[3][16][30] , \s_mux2_signals[3][16][29] , 
        \s_mux2_signals[3][16][28] , \s_mux2_signals[3][16][27] , 
        \s_mux2_signals[3][16][26] , \s_mux2_signals[3][16][25] , 
        \s_mux2_signals[3][16][24] , \s_mux2_signals[3][16][23] , 
        \s_mux2_signals[3][16][22] , \s_mux2_signals[3][16][21] , 
        \s_mux2_signals[3][16][20] , \s_mux2_signals[3][16][19] , 
        \s_mux2_signals[3][16][18] , \s_mux2_signals[3][16][17] , 
        \s_mux2_signals[3][16][16] , \s_mux2_signals[3][16][15] , 
        \s_mux2_signals[3][16][14] , \s_mux2_signals[3][16][13] , 
        \s_mux2_signals[3][16][12] , \s_mux2_signals[3][16][11] , 
        \s_mux2_signals[3][16][10] , \s_mux2_signals[3][16][9] , 
        \s_mux2_signals[3][16][8] , \s_mux2_signals[3][16][7] , 
        \s_mux2_signals[3][16][6] , \s_mux2_signals[3][16][5] , 
        \s_mux2_signals[3][16][4] , \s_mux2_signals[3][16][3] , 
        \s_mux2_signals[3][16][2] , \s_mux2_signals[3][16][1] , 
        \s_mux2_signals[3][16][0] }), .port1({\s_mux2_signals[3][24][31] , 
        \s_mux2_signals[3][24][30] , \s_mux2_signals[3][24][29] , 
        \s_mux2_signals[3][24][28] , \s_mux2_signals[3][24][27] , 
        \s_mux2_signals[3][24][26] , \s_mux2_signals[3][24][25] , 
        \s_mux2_signals[3][24][24] , \s_mux2_signals[3][24][23] , 
        \s_mux2_signals[3][24][22] , \s_mux2_signals[3][24][21] , 
        \s_mux2_signals[3][24][20] , \s_mux2_signals[3][24][19] , 
        \s_mux2_signals[3][24][18] , \s_mux2_signals[3][24][17] , 
        \s_mux2_signals[3][24][16] , \s_mux2_signals[3][24][15] , 
        \s_mux2_signals[3][24][14] , \s_mux2_signals[3][24][13] , 
        \s_mux2_signals[3][24][12] , \s_mux2_signals[3][24][11] , 
        \s_mux2_signals[3][24][10] , \s_mux2_signals[3][24][9] , 
        \s_mux2_signals[3][24][8] , \s_mux2_signals[3][24][7] , 
        \s_mux2_signals[3][24][6] , \s_mux2_signals[3][24][5] , 
        \s_mux2_signals[3][24][4] , \s_mux2_signals[3][24][3] , 
        \s_mux2_signals[3][24][2] , \s_mux2_signals[3][24][1] , 
        \s_mux2_signals[3][24][0] }), .sel(s_addrRd2_Fei_Tmux[3]), .portY({
        \s_mux2_signals[4][16][31] , \s_mux2_signals[4][16][30] , 
        \s_mux2_signals[4][16][29] , \s_mux2_signals[4][16][28] , 
        \s_mux2_signals[4][16][27] , \s_mux2_signals[4][16][26] , 
        \s_mux2_signals[4][16][25] , \s_mux2_signals[4][16][24] , 
        \s_mux2_signals[4][16][23] , \s_mux2_signals[4][16][22] , 
        \s_mux2_signals[4][16][21] , \s_mux2_signals[4][16][20] , 
        \s_mux2_signals[4][16][19] , \s_mux2_signals[4][16][18] , 
        \s_mux2_signals[4][16][17] , \s_mux2_signals[4][16][16] , 
        \s_mux2_signals[4][16][15] , \s_mux2_signals[4][16][14] , 
        \s_mux2_signals[4][16][13] , \s_mux2_signals[4][16][12] , 
        \s_mux2_signals[4][16][11] , \s_mux2_signals[4][16][10] , 
        \s_mux2_signals[4][16][9] , \s_mux2_signals[4][16][8] , 
        \s_mux2_signals[4][16][7] , \s_mux2_signals[4][16][6] , 
        \s_mux2_signals[4][16][5] , \s_mux2_signals[4][16][4] , 
        \s_mux2_signals[4][16][3] , \s_mux2_signals[4][16][2] , 
        \s_mux2_signals[4][16][1] , \s_mux2_signals[4][16][0] }) );
  Mux_NBit_2x1_NBIT_IN32_18 MUX2_4_0 ( .port0({\s_mux2_signals[4][0][31] , 
        \s_mux2_signals[4][0][30] , \s_mux2_signals[4][0][29] , 
        \s_mux2_signals[4][0][28] , \s_mux2_signals[4][0][27] , 
        \s_mux2_signals[4][0][26] , \s_mux2_signals[4][0][25] , 
        \s_mux2_signals[4][0][24] , \s_mux2_signals[4][0][23] , 
        \s_mux2_signals[4][0][22] , \s_mux2_signals[4][0][21] , 
        \s_mux2_signals[4][0][20] , \s_mux2_signals[4][0][19] , 
        \s_mux2_signals[4][0][18] , \s_mux2_signals[4][0][17] , 
        \s_mux2_signals[4][0][16] , \s_mux2_signals[4][0][15] , 
        \s_mux2_signals[4][0][14] , \s_mux2_signals[4][0][13] , 
        \s_mux2_signals[4][0][12] , \s_mux2_signals[4][0][11] , 
        \s_mux2_signals[4][0][10] , \s_mux2_signals[4][0][9] , 
        \s_mux2_signals[4][0][8] , \s_mux2_signals[4][0][7] , 
        \s_mux2_signals[4][0][6] , \s_mux2_signals[4][0][5] , 
        \s_mux2_signals[4][0][4] , \s_mux2_signals[4][0][3] , 
        \s_mux2_signals[4][0][2] , \s_mux2_signals[4][0][1] , 
        \s_mux2_signals[4][0][0] }), .port1({\s_mux2_signals[4][16][31] , 
        \s_mux2_signals[4][16][30] , \s_mux2_signals[4][16][29] , 
        \s_mux2_signals[4][16][28] , \s_mux2_signals[4][16][27] , 
        \s_mux2_signals[4][16][26] , \s_mux2_signals[4][16][25] , 
        \s_mux2_signals[4][16][24] , \s_mux2_signals[4][16][23] , 
        \s_mux2_signals[4][16][22] , \s_mux2_signals[4][16][21] , 
        \s_mux2_signals[4][16][20] , \s_mux2_signals[4][16][19] , 
        \s_mux2_signals[4][16][18] , \s_mux2_signals[4][16][17] , 
        \s_mux2_signals[4][16][16] , \s_mux2_signals[4][16][15] , 
        \s_mux2_signals[4][16][14] , \s_mux2_signals[4][16][13] , 
        \s_mux2_signals[4][16][12] , \s_mux2_signals[4][16][11] , 
        \s_mux2_signals[4][16][10] , \s_mux2_signals[4][16][9] , 
        \s_mux2_signals[4][16][8] , \s_mux2_signals[4][16][7] , 
        \s_mux2_signals[4][16][6] , \s_mux2_signals[4][16][5] , 
        \s_mux2_signals[4][16][4] , \s_mux2_signals[4][16][3] , 
        \s_mux2_signals[4][16][2] , \s_mux2_signals[4][16][1] , 
        \s_mux2_signals[4][16][0] }), .sel(s_addrRd2_Fei_Tmux[4]), .portY(
        RF_out2) );
  CLKBUF_X1 U2 ( .A(\s_mux2_signals[0][31][0] ), .Z(n21) );
  CLKBUF_X1 U3 ( .A(RF_data_in[27]), .Z(n109) );
  CLKBUF_X1 U4 ( .A(RF_data_in[28]), .Z(n110) );
  CLKBUF_X1 U6 ( .A(RF_data_in[29]), .Z(n111) );
  BUF_X1 U7 ( .A(RF_reset), .Z(n117) );
  BUF_X1 U8 ( .A(RF_reset), .Z(n118) );
  CLKBUF_X1 U9 ( .A(RF_data_in[19]), .Z(n89) );
  CLKBUF_X1 U10 ( .A(RF_data_in[20]), .Z(n92) );
  CLKBUF_X1 U11 ( .A(RF_data_in[21]), .Z(n95) );
  CLKBUF_X1 U12 ( .A(RF_data_in[23]), .Z(n99) );
  CLKBUF_X1 U13 ( .A(RF_data_in[24]), .Z(n102) );
  CLKBUF_X1 U14 ( .A(RF_data_in[25]), .Z(n105) );
  CLKBUF_X1 U15 ( .A(RF_data_in[19]), .Z(n90) );
  CLKBUF_X1 U16 ( .A(RF_data_in[20]), .Z(n93) );
  CLKBUF_X1 U17 ( .A(RF_data_in[21]), .Z(n96) );
  CLKBUF_X1 U18 ( .A(RF_data_in[23]), .Z(n100) );
  CLKBUF_X1 U19 ( .A(RF_data_in[24]), .Z(n103) );
  CLKBUF_X1 U20 ( .A(RF_data_in[25]), .Z(n106) );
  CLKBUF_X1 U21 ( .A(RF_data_in[1]), .Z(n37) );
  CLKBUF_X1 U22 ( .A(RF_data_in[19]), .Z(n91) );
  CLKBUF_X1 U23 ( .A(RF_data_in[20]), .Z(n94) );
  CLKBUF_X1 U24 ( .A(RF_data_in[21]), .Z(n97) );
  CLKBUF_X1 U25 ( .A(RF_data_in[22]), .Z(n98) );
  CLKBUF_X1 U26 ( .A(RF_data_in[23]), .Z(n101) );
  CLKBUF_X1 U27 ( .A(RF_data_in[24]), .Z(n104) );
  CLKBUF_X1 U28 ( .A(RF_data_in[25]), .Z(n107) );
  CLKBUF_X1 U29 ( .A(RF_data_in[26]), .Z(n108) );
  CLKBUF_X1 U30 ( .A(RF_data_in[7]), .Z(n53) );
  CLKBUF_X1 U31 ( .A(RF_data_in[7]), .Z(n54) );
  CLKBUF_X1 U32 ( .A(RF_data_in[7]), .Z(n55) );
  BUF_X1 U33 ( .A(RF_reset), .Z(n119) );
  CLKBUF_X1 U34 ( .A(RF_data_in[2]), .Z(n38) );
  CLKBUF_X1 U35 ( .A(RF_data_in[3]), .Z(n41) );
  CLKBUF_X1 U36 ( .A(RF_data_in[4]), .Z(n44) );
  CLKBUF_X1 U37 ( .A(RF_data_in[5]), .Z(n47) );
  CLKBUF_X1 U38 ( .A(RF_data_in[6]), .Z(n50) );
  CLKBUF_X1 U39 ( .A(RF_data_in[8]), .Z(n56) );
  CLKBUF_X1 U40 ( .A(RF_data_in[9]), .Z(n59) );
  CLKBUF_X1 U41 ( .A(RF_data_in[10]), .Z(n62) );
  CLKBUF_X1 U42 ( .A(RF_data_in[11]), .Z(n65) );
  CLKBUF_X1 U43 ( .A(RF_data_in[12]), .Z(n68) );
  CLKBUF_X1 U44 ( .A(RF_data_in[13]), .Z(n71) );
  CLKBUF_X1 U45 ( .A(RF_data_in[14]), .Z(n74) );
  CLKBUF_X1 U46 ( .A(RF_data_in[15]), .Z(n77) );
  CLKBUF_X1 U47 ( .A(RF_data_in[16]), .Z(n80) );
  CLKBUF_X1 U48 ( .A(RF_data_in[17]), .Z(n83) );
  CLKBUF_X1 U49 ( .A(RF_data_in[18]), .Z(n86) );
  CLKBUF_X1 U50 ( .A(RF_data_in[2]), .Z(n39) );
  CLKBUF_X1 U51 ( .A(RF_data_in[3]), .Z(n42) );
  CLKBUF_X1 U52 ( .A(RF_data_in[4]), .Z(n45) );
  CLKBUF_X1 U53 ( .A(RF_data_in[5]), .Z(n48) );
  CLKBUF_X1 U54 ( .A(RF_data_in[6]), .Z(n51) );
  CLKBUF_X1 U55 ( .A(RF_data_in[8]), .Z(n57) );
  CLKBUF_X1 U56 ( .A(RF_data_in[9]), .Z(n60) );
  CLKBUF_X1 U57 ( .A(RF_data_in[10]), .Z(n63) );
  CLKBUF_X1 U58 ( .A(RF_data_in[11]), .Z(n66) );
  CLKBUF_X1 U59 ( .A(RF_data_in[12]), .Z(n69) );
  CLKBUF_X1 U60 ( .A(RF_data_in[13]), .Z(n72) );
  CLKBUF_X1 U61 ( .A(RF_data_in[14]), .Z(n75) );
  CLKBUF_X1 U62 ( .A(RF_data_in[15]), .Z(n78) );
  CLKBUF_X1 U63 ( .A(RF_data_in[16]), .Z(n81) );
  CLKBUF_X1 U64 ( .A(RF_data_in[17]), .Z(n84) );
  CLKBUF_X1 U65 ( .A(RF_data_in[18]), .Z(n87) );
  CLKBUF_X1 U66 ( .A(RF_data_in[30]), .Z(n112) );
  CLKBUF_X1 U67 ( .A(RF_data_in[0]), .Z(n36) );
  CLKBUF_X1 U68 ( .A(RF_data_in[2]), .Z(n40) );
  CLKBUF_X1 U69 ( .A(RF_data_in[3]), .Z(n43) );
  CLKBUF_X1 U70 ( .A(RF_data_in[4]), .Z(n46) );
  CLKBUF_X1 U71 ( .A(RF_data_in[5]), .Z(n49) );
  CLKBUF_X1 U72 ( .A(RF_data_in[6]), .Z(n52) );
  CLKBUF_X1 U73 ( .A(RF_data_in[8]), .Z(n58) );
  CLKBUF_X1 U74 ( .A(RF_data_in[9]), .Z(n61) );
  CLKBUF_X1 U75 ( .A(RF_data_in[10]), .Z(n64) );
  CLKBUF_X1 U76 ( .A(RF_data_in[11]), .Z(n67) );
  CLKBUF_X1 U77 ( .A(RF_data_in[12]), .Z(n70) );
  CLKBUF_X1 U78 ( .A(RF_data_in[13]), .Z(n73) );
  CLKBUF_X1 U79 ( .A(RF_data_in[14]), .Z(n76) );
  CLKBUF_X1 U80 ( .A(RF_data_in[15]), .Z(n79) );
  CLKBUF_X1 U81 ( .A(RF_data_in[16]), .Z(n82) );
  CLKBUF_X1 U82 ( .A(RF_data_in[17]), .Z(n85) );
  CLKBUF_X1 U83 ( .A(RF_data_in[18]), .Z(n88) );
  BUF_X1 U84 ( .A(n4), .Z(n22) );
  BUF_X1 U85 ( .A(n4), .Z(n23) );
  CLKBUF_X1 U86 ( .A(RF_enable), .Z(n116) );
  BUF_X1 U87 ( .A(n4), .Z(n24) );
  BUF_X1 U88 ( .A(n2), .Z(n26) );
  BUF_X1 U89 ( .A(n2), .Z(n25) );
  BUF_X1 U90 ( .A(n2), .Z(n27) );
  CLKBUF_X1 U91 ( .A(RF_enable), .Z(n114) );
  CLKBUF_X1 U92 ( .A(RF_enable), .Z(n115) );
  AND2_X1 U93 ( .A1(RF_RD1), .A2(n116), .ZN(s_rd1_enable) );
  BUF_X1 U94 ( .A(s_addrRd1_Fei_Tmux[2]), .Z(n35) );
  AND2_X1 U95 ( .A1(n116), .A2(RF_WR), .ZN(s_wr_enable) );
  AND2_X1 U96 ( .A1(RF_RD2), .A2(n116), .ZN(s_rd2_enable) );
  BUF_X1 U97 ( .A(s_addrRd2_Fei_Tmux[2]), .Z(n31) );
  CLKBUF_X1 U98 ( .A(RF_data_in[31]), .Z(n113) );
  CLKBUF_X1 U99 ( .A(s_addrRd2_Fei_Tmux[1]), .Z(n28) );
  CLKBUF_X1 U100 ( .A(s_addrRd2_Fei_Tmux[1]), .Z(n29) );
  CLKBUF_X1 U101 ( .A(s_addrRd2_Fei_Tmux[1]), .Z(n30) );
  CLKBUF_X1 U102 ( .A(s_addrRd1_Fei_Tmux[1]), .Z(n32) );
  CLKBUF_X1 U103 ( .A(s_addrRd1_Fei_Tmux[1]), .Z(n33) );
  CLKBUF_X1 U104 ( .A(s_addrRd1_Fei_Tmux[1]), .Z(n34) );
endmodule


module NRegister_N5_3 ( clk, reset, data_in, enable, load, data_out );
  input [4:0] data_in;
  output [4:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, net110627, net110628, net110629, net110630,
         net110631, n14, n15, n16, n17, n18, n19, n20, n8;

  DFFR_X1 \data_out_reg[4]  ( .D(n2), .CK(clk), .RN(n8), .Q(data_out[4]), .QN(
        net110631) );
  DFFR_X1 \data_out_reg[3]  ( .D(n4), .CK(clk), .RN(n8), .Q(data_out[3]), .QN(
        net110630) );
  DFFR_X1 \data_out_reg[2]  ( .D(n5), .CK(clk), .RN(n8), .Q(data_out[2]), .QN(
        net110629) );
  DFFR_X1 \data_out_reg[1]  ( .D(n6), .CK(clk), .RN(n8), .Q(data_out[1]), .QN(
        net110628) );
  DFFR_X1 \data_out_reg[0]  ( .D(n7), .CK(clk), .RN(n8), .Q(data_out[0]), .QN(
        net110627) );
  INV_X1 U3 ( .A(n14), .ZN(n16) );
  NAND2_X1 U4 ( .A1(load), .A2(enable), .ZN(n14) );
  OAI22_X1 U5 ( .A1(n14), .A2(n15), .B1(net110627), .B2(n16), .ZN(n7) );
  INV_X1 U6 ( .A(data_in[0]), .ZN(n15) );
  OAI22_X1 U7 ( .A1(n14), .A2(n17), .B1(net110628), .B2(n16), .ZN(n6) );
  INV_X1 U8 ( .A(data_in[1]), .ZN(n17) );
  OAI22_X1 U9 ( .A1(n14), .A2(n18), .B1(net110629), .B2(n16), .ZN(n5) );
  INV_X1 U10 ( .A(data_in[2]), .ZN(n18) );
  OAI22_X1 U11 ( .A1(n14), .A2(n19), .B1(net110630), .B2(n16), .ZN(n4) );
  INV_X1 U12 ( .A(data_in[3]), .ZN(n19) );
  OAI22_X1 U13 ( .A1(n14), .A2(n20), .B1(net110631), .B2(n16), .ZN(n2) );
  INV_X1 U14 ( .A(data_in[4]), .ZN(n20) );
  INV_X1 U15 ( .A(reset), .ZN(n8) );
endmodule


module NRegister_N5_0 ( clk, reset, data_in, enable, load, data_out );
  input [4:0] data_in;
  output [4:0] data_out;
  input clk, reset, enable, load;
  wire   n14, n15, n16, n17, n19, net106790, net106791, net106792, net106793,
         net106794, n8, n9, n10, n11, n12, n13, n20, n2;

  DFFR_X1 \data_out_reg[4]  ( .D(n19), .CK(clk), .RN(n2), .Q(data_out[4]), 
        .QN(net106794) );
  DFFR_X1 \data_out_reg[3]  ( .D(n17), .CK(clk), .RN(n2), .Q(data_out[3]), 
        .QN(net106793) );
  DFFR_X1 \data_out_reg[2]  ( .D(n16), .CK(clk), .RN(n2), .Q(data_out[2]), 
        .QN(net106792) );
  DFFR_X1 \data_out_reg[1]  ( .D(n15), .CK(clk), .RN(n2), .Q(data_out[1]), 
        .QN(net106791) );
  DFFR_X1 \data_out_reg[0]  ( .D(n14), .CK(clk), .RN(n2), .Q(data_out[0]), 
        .QN(net106790) );
  INV_X1 U3 ( .A(n8), .ZN(n10) );
  NAND2_X1 U4 ( .A1(load), .A2(enable), .ZN(n8) );
  OAI22_X1 U5 ( .A1(n8), .A2(n20), .B1(net106790), .B2(n10), .ZN(n14) );
  INV_X1 U6 ( .A(data_in[0]), .ZN(n20) );
  OAI22_X1 U7 ( .A1(n8), .A2(n13), .B1(net106791), .B2(n10), .ZN(n15) );
  INV_X1 U8 ( .A(data_in[1]), .ZN(n13) );
  OAI22_X1 U9 ( .A1(n8), .A2(n12), .B1(net106792), .B2(n10), .ZN(n16) );
  INV_X1 U10 ( .A(data_in[2]), .ZN(n12) );
  OAI22_X1 U11 ( .A1(n8), .A2(n11), .B1(net106793), .B2(n10), .ZN(n17) );
  INV_X1 U12 ( .A(data_in[3]), .ZN(n11) );
  OAI22_X1 U13 ( .A1(n8), .A2(n9), .B1(net106794), .B2(n10), .ZN(n19) );
  INV_X1 U14 ( .A(data_in[4]), .ZN(n9) );
  INV_X1 U15 ( .A(reset), .ZN(n2) );
endmodule


module PropagateCarryLookahead_N32_0 ( A, B, Cin, Sum, Cout );
  input [31:0] A;
  input [31:0] B;
  output [31:0] Sum;
  input Cin;
  output Cout;

  wire   [31:0] s_G1;
  wire   [31:0] s_P1;
  wire   [31:0] s_G2;
  wire   [31:0] s_P2;
  wire   SYNOPSYS_UNCONNECTED__0;

  PG_network_N32_0 PG ( .A(A), .B(B), .c_in(1'b0), .G(s_G1), .P({s_P1[31:1], 
        SYNOPSYS_UNCONNECTED__0}) );
  Carry_Network_N32_0 CN ( .G(s_G1), .P({s_P1[31:1], 1'b0}), .Cin(Cin), .Cout(
        Cout), .Gout(s_G2), .Pout(s_P2) );
  Sum_Network_N32_0 SN ( .G(s_G2), .P(s_P2), .S(Sum) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_121 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n4, n5, n6, n7, n8, n9, n10, n11,
         n12, n13, n14, n15, n16, n17;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n17), .ZN(n7) );
  INV_X1 U2 ( .A(n17), .ZN(n8) );
  BUF_X1 U3 ( .A(n4), .Z(n9) );
  BUF_X1 U4 ( .A(n6), .Z(n15) );
  BUF_X1 U5 ( .A(n5), .Z(n14) );
  BUF_X1 U6 ( .A(n5), .Z(n12) );
  BUF_X1 U7 ( .A(n4), .Z(n11) );
  BUF_X1 U8 ( .A(n5), .Z(n13) );
  BUF_X1 U9 ( .A(n4), .Z(n10) );
  BUF_X1 U10 ( .A(n6), .Z(n17) );
  BUF_X1 U11 ( .A(n6), .Z(n16) );
  INV_X1 U12 ( .A(n34), .ZN(N9) );
  INV_X1 U13 ( .A(n40), .ZN(N4) );
  INV_X1 U14 ( .A(n39), .ZN(N5) );
  INV_X1 U15 ( .A(n38), .ZN(N6) );
  INV_X1 U16 ( .A(n37), .ZN(N7) );
  INV_X1 U17 ( .A(n36), .ZN(N8) );
  INV_X1 U18 ( .A(n42), .ZN(N32) );
  INV_X1 U19 ( .A(n41), .ZN(N33) );
  BUF_X1 U20 ( .A(sel), .Z(n6) );
  BUF_X1 U21 ( .A(sel), .Z(n5) );
  BUF_X1 U22 ( .A(sel), .Z(n4) );
  INV_X1 U23 ( .A(n56), .ZN(N2) );
  INV_X1 U24 ( .A(n45), .ZN(N3) );
  INV_X1 U25 ( .A(n63), .ZN(N13) );
  INV_X1 U26 ( .A(n62), .ZN(N14) );
  INV_X1 U27 ( .A(n61), .ZN(N15) );
  INV_X1 U28 ( .A(n60), .ZN(N16) );
  INV_X1 U29 ( .A(n59), .ZN(N17) );
  INV_X1 U30 ( .A(n58), .ZN(N18) );
  INV_X1 U31 ( .A(n57), .ZN(N19) );
  INV_X1 U32 ( .A(n55), .ZN(N20) );
  INV_X1 U33 ( .A(n54), .ZN(N21) );
  INV_X1 U34 ( .A(n53), .ZN(N22) );
  INV_X1 U35 ( .A(n52), .ZN(N23) );
  INV_X1 U36 ( .A(n51), .ZN(N24) );
  INV_X1 U37 ( .A(n50), .ZN(N25) );
  INV_X1 U38 ( .A(n49), .ZN(N26) );
  INV_X1 U39 ( .A(n48), .ZN(N27) );
  INV_X1 U40 ( .A(n47), .ZN(N28) );
  INV_X1 U41 ( .A(n46), .ZN(N29) );
  INV_X1 U42 ( .A(n44), .ZN(N30) );
  INV_X1 U43 ( .A(n43), .ZN(N31) );
  INV_X1 U44 ( .A(n66), .ZN(N10) );
  INV_X1 U45 ( .A(n65), .ZN(N11) );
  INV_X1 U46 ( .A(n64), .ZN(N12) );
  AOI22_X1 U47 ( .A1(port0[2]), .A2(n7), .B1(port1[2]), .B2(n10), .ZN(n40) );
  AOI22_X1 U48 ( .A1(port0[3]), .A2(n8), .B1(port1[3]), .B2(n9), .ZN(n39) );
  AOI22_X1 U49 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(n9), .ZN(n38) );
  AOI22_X1 U50 ( .A1(port0[5]), .A2(n8), .B1(port1[5]), .B2(n9), .ZN(n37) );
  AOI22_X1 U51 ( .A1(port0[6]), .A2(n8), .B1(port1[6]), .B2(n9), .ZN(n36) );
  AOI22_X1 U52 ( .A1(port0[7]), .A2(n7), .B1(n16), .B2(port1[7]), .ZN(n34) );
  AOI22_X1 U53 ( .A1(port0[30]), .A2(n8), .B1(port1[30]), .B2(n10), .ZN(n42)
         );
  AOI22_X1 U54 ( .A1(port0[31]), .A2(n7), .B1(port1[31]), .B2(n10), .ZN(n41)
         );
  AOI22_X1 U55 ( .A1(port0[0]), .A2(n7), .B1(port1[0]), .B2(n14), .ZN(n56) );
  AOI22_X1 U56 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(n11), .ZN(n45) );
  AOI22_X1 U57 ( .A1(port0[8]), .A2(n7), .B1(port1[8]), .B2(n16), .ZN(n66) );
  AOI22_X1 U58 ( .A1(port0[9]), .A2(n7), .B1(port1[9]), .B2(n16), .ZN(n65) );
  AOI22_X1 U59 ( .A1(port0[10]), .A2(n7), .B1(port1[10]), .B2(n16), .ZN(n64)
         );
  AOI22_X1 U60 ( .A1(port0[11]), .A2(n7), .B1(port1[11]), .B2(n15), .ZN(n63)
         );
  AOI22_X1 U61 ( .A1(port0[12]), .A2(n7), .B1(port1[12]), .B2(n15), .ZN(n62)
         );
  AOI22_X1 U62 ( .A1(port0[13]), .A2(n7), .B1(port1[13]), .B2(n15), .ZN(n61)
         );
  AOI22_X1 U63 ( .A1(port0[14]), .A2(n7), .B1(port1[14]), .B2(n15), .ZN(n60)
         );
  AOI22_X1 U64 ( .A1(port0[15]), .A2(n7), .B1(port1[15]), .B2(n14), .ZN(n59)
         );
  AOI22_X1 U65 ( .A1(port0[16]), .A2(n7), .B1(port1[16]), .B2(n14), .ZN(n58)
         );
  AOI22_X1 U66 ( .A1(port0[17]), .A2(n7), .B1(port1[17]), .B2(n14), .ZN(n57)
         );
  AOI22_X1 U67 ( .A1(port0[18]), .A2(n7), .B1(port1[18]), .B2(n13), .ZN(n55)
         );
  AOI22_X1 U68 ( .A1(port0[19]), .A2(n8), .B1(port1[19]), .B2(n13), .ZN(n54)
         );
  AOI22_X1 U69 ( .A1(port0[20]), .A2(n8), .B1(port1[20]), .B2(n13), .ZN(n53)
         );
  AOI22_X1 U70 ( .A1(port0[21]), .A2(n8), .B1(port1[21]), .B2(n12), .ZN(n52)
         );
  AOI22_X1 U71 ( .A1(port0[22]), .A2(n8), .B1(port1[22]), .B2(n12), .ZN(n51)
         );
  AOI22_X1 U72 ( .A1(port0[23]), .A2(n8), .B1(port1[23]), .B2(n12), .ZN(n50)
         );
  AOI22_X1 U73 ( .A1(port0[24]), .A2(n8), .B1(port1[24]), .B2(n12), .ZN(n49)
         );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n8), .B1(port1[25]), .B2(n11), .ZN(n48)
         );
  AOI22_X1 U75 ( .A1(port0[26]), .A2(n8), .B1(port1[26]), .B2(n11), .ZN(n47)
         );
  AOI22_X1 U76 ( .A1(port0[27]), .A2(n8), .B1(port1[27]), .B2(n11), .ZN(n46)
         );
  AOI22_X1 U77 ( .A1(port0[28]), .A2(n8), .B1(port1[28]), .B2(n10), .ZN(n44)
         );
  AOI22_X1 U78 ( .A1(port0[29]), .A2(n8), .B1(port1[29]), .B2(n13), .ZN(n43)
         );
endmodule


module Mux_1Bit_2X1_4 ( port0, port1, sel, portY );
  input port0, port1, sel;
  output portY;
  wire   n3, n4;

  INV_X4 U1 ( .A(n3), .ZN(portY) );
  AOI22_X1 U2 ( .A1(port0), .A2(n4), .B1(sel), .B2(port1), .ZN(n3) );
  INV_X1 U3 ( .A(sel), .ZN(n4) );
endmodule


module Mux_Bit_NBIT_Sel5 ( inputs, sel, \output  );
  input [31:0] inputs;
  input [4:0] sel;
  output \output ;
  wire   n14, n16, n17, n18, n20, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55;

  NOR2_X1 U1 ( .A1(n52), .A2(n51), .ZN(n24) );
  NOR2_X1 U2 ( .A1(n51), .A2(sel[1]), .ZN(n28) );
  NOR2_X1 U3 ( .A1(sel[0]), .A2(sel[1]), .ZN(n27) );
  NOR2_X1 U4 ( .A1(n52), .A2(sel[0]), .ZN(n23) );
  INV_X1 U5 ( .A(sel[1]), .ZN(n52) );
  AOI221_X1 U6 ( .B1(inputs[2]), .B2(n23), .C1(inputs[3]), .C2(n24), .A(n25), 
        .ZN(n22) );
  INV_X1 U7 ( .A(n26), .ZN(n25) );
  AOI22_X1 U8 ( .A1(inputs[0]), .A2(n27), .B1(inputs[1]), .B2(n28), .ZN(n26)
         );
  AOI221_X1 U9 ( .B1(inputs[10]), .B2(n23), .C1(inputs[11]), .C2(n24), .A(n33), 
        .ZN(n32) );
  INV_X1 U10 ( .A(n34), .ZN(n33) );
  AOI22_X1 U11 ( .A1(inputs[8]), .A2(n27), .B1(inputs[9]), .B2(n28), .ZN(n34)
         );
  AOI221_X1 U12 ( .B1(inputs[18]), .B2(n23), .C1(inputs[19]), .C2(n24), .A(n41), .ZN(n40) );
  INV_X1 U13 ( .A(n42), .ZN(n41) );
  AOI22_X1 U14 ( .A1(inputs[16]), .A2(n27), .B1(inputs[17]), .B2(n28), .ZN(n42) );
  AOI221_X1 U15 ( .B1(inputs[26]), .B2(n23), .C1(inputs[27]), .C2(n24), .A(n47), .ZN(n46) );
  INV_X1 U16 ( .A(n48), .ZN(n47) );
  AOI22_X1 U17 ( .A1(inputs[24]), .A2(n27), .B1(inputs[25]), .B2(n28), .ZN(n48) );
  AOI221_X1 U18 ( .B1(inputs[6]), .B2(n23), .C1(inputs[7]), .C2(n24), .A(n29), 
        .ZN(n20) );
  INV_X1 U19 ( .A(n30), .ZN(n29) );
  AOI22_X1 U20 ( .A1(inputs[4]), .A2(n27), .B1(inputs[5]), .B2(n28), .ZN(n30)
         );
  AOI221_X1 U21 ( .B1(inputs[22]), .B2(n23), .C1(inputs[23]), .C2(n24), .A(n43), .ZN(n39) );
  INV_X1 U22 ( .A(n44), .ZN(n43) );
  AOI22_X1 U23 ( .A1(inputs[20]), .A2(n27), .B1(inputs[21]), .B2(n28), .ZN(n44) );
  AOI22_X1 U24 ( .A1(sel[3]), .A2(n17), .B1(n18), .B2(n54), .ZN(n16) );
  OAI22_X1 U25 ( .A1(n31), .A2(n53), .B1(sel[2]), .B2(n32), .ZN(n17) );
  OAI22_X1 U26 ( .A1(n20), .A2(n53), .B1(sel[2]), .B2(n22), .ZN(n18) );
  AOI221_X1 U27 ( .B1(inputs[14]), .B2(n23), .C1(inputs[15]), .C2(n24), .A(n35), .ZN(n31) );
  OAI22_X1 U28 ( .A1(n14), .A2(n55), .B1(sel[4]), .B2(n16), .ZN(\output ) );
  AOI22_X1 U29 ( .A1(sel[3]), .A2(n37), .B1(n38), .B2(n54), .ZN(n14) );
  OAI22_X1 U30 ( .A1(n45), .A2(n53), .B1(sel[2]), .B2(n46), .ZN(n37) );
  OAI22_X1 U31 ( .A1(n39), .A2(n53), .B1(sel[2]), .B2(n40), .ZN(n38) );
  AOI221_X1 U32 ( .B1(inputs[30]), .B2(n23), .C1(inputs[31]), .C2(n24), .A(n49), .ZN(n45) );
  INV_X1 U33 ( .A(n36), .ZN(n35) );
  AOI22_X1 U34 ( .A1(inputs[12]), .A2(n27), .B1(inputs[13]), .B2(n28), .ZN(n36) );
  INV_X1 U35 ( .A(n50), .ZN(n49) );
  AOI22_X1 U36 ( .A1(inputs[28]), .A2(n27), .B1(inputs[29]), .B2(n28), .ZN(n50) );
  INV_X1 U37 ( .A(sel[0]), .ZN(n51) );
  INV_X1 U38 ( .A(sel[2]), .ZN(n53) );
  INV_X1 U39 ( .A(sel[3]), .ZN(n54) );
  INV_X1 U40 ( .A(sel[4]), .ZN(n55) );
endmodule


module SAT_Counter_BTB_N3_0 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, 
        SAT_update, SAT_setToDef, SAT_SO );
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  output SAT_SO;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;
  wire   [1:0] s_cnt;

  UD_COUNTER_BTB_UDC_NBIT3_0 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), .UDC_CLK(
        s_clk), .UDC_RST(s_reset), .UDC_OUT({SAT_SO, s_cnt}) );
  CU_SatCounter_32 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  AND3_X1 U1 ( .A1(s_cnt[1]), .A2(SAT_SO), .A3(s_cnt[0]), .ZN(s_TcMax) );
  NOR3_X1 U2 ( .A1(SAT_SO), .A2(s_cnt[1]), .A3(s_cnt[0]), .ZN(s_TcMin) );
endmodule


module NRotateRegister_N32 ( clk, reset, enable, load, data_in, rotate, 
        data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load, rotate;
  wire   n2, n3, n4, n5, n6, n7, n8;
  wire   [1:0] s_phi;
  wire   [31:0] s_D_Fmux_TFF;

  D_FF_0 DFF_i_0 ( .D(s_D_Fmux_TFF[0]), .clk(clk), .Q(data_out[0]) );
  D_FF_31 DFF_i_1 ( .D(s_D_Fmux_TFF[1]), .clk(clk), .Q(data_out[1]) );
  D_FF_30 DFF_i_2 ( .D(s_D_Fmux_TFF[2]), .clk(clk), .Q(data_out[2]) );
  D_FF_29 DFF_i_3 ( .D(s_D_Fmux_TFF[3]), .clk(clk), .Q(data_out[3]) );
  D_FF_28 DFF_i_4 ( .D(s_D_Fmux_TFF[4]), .clk(clk), .Q(data_out[4]) );
  D_FF_27 DFF_i_5 ( .D(s_D_Fmux_TFF[5]), .clk(clk), .Q(data_out[5]) );
  D_FF_26 DFF_i_6 ( .D(s_D_Fmux_TFF[6]), .clk(clk), .Q(data_out[6]) );
  D_FF_25 DFF_i_7 ( .D(s_D_Fmux_TFF[7]), .clk(clk), .Q(data_out[7]) );
  D_FF_24 DFF_i_8 ( .D(s_D_Fmux_TFF[8]), .clk(clk), .Q(data_out[8]) );
  D_FF_23 DFF_i_9 ( .D(s_D_Fmux_TFF[9]), .clk(clk), .Q(data_out[9]) );
  D_FF_22 DFF_i_10 ( .D(s_D_Fmux_TFF[10]), .clk(clk), .Q(data_out[10]) );
  D_FF_21 DFF_i_11 ( .D(s_D_Fmux_TFF[11]), .clk(clk), .Q(data_out[11]) );
  D_FF_20 DFF_i_12 ( .D(s_D_Fmux_TFF[12]), .clk(clk), .Q(data_out[12]) );
  D_FF_19 DFF_i_13 ( .D(s_D_Fmux_TFF[13]), .clk(clk), .Q(data_out[13]) );
  D_FF_18 DFF_i_14 ( .D(s_D_Fmux_TFF[14]), .clk(clk), .Q(data_out[14]) );
  D_FF_17 DFF_i_15 ( .D(s_D_Fmux_TFF[15]), .clk(clk), .Q(data_out[15]) );
  D_FF_16 DFF_i_16 ( .D(s_D_Fmux_TFF[16]), .clk(clk), .Q(data_out[16]) );
  D_FF_15 DFF_i_17 ( .D(s_D_Fmux_TFF[17]), .clk(clk), .Q(data_out[17]) );
  D_FF_14 DFF_i_18 ( .D(s_D_Fmux_TFF[18]), .clk(clk), .Q(data_out[18]) );
  D_FF_13 DFF_i_19 ( .D(s_D_Fmux_TFF[19]), .clk(clk), .Q(data_out[19]) );
  D_FF_12 DFF_i_20 ( .D(s_D_Fmux_TFF[20]), .clk(clk), .Q(data_out[20]) );
  D_FF_11 DFF_i_21 ( .D(s_D_Fmux_TFF[21]), .clk(clk), .Q(data_out[21]) );
  D_FF_10 DFF_i_22 ( .D(s_D_Fmux_TFF[22]), .clk(clk), .Q(data_out[22]) );
  D_FF_9 DFF_i_23 ( .D(s_D_Fmux_TFF[23]), .clk(clk), .Q(data_out[23]) );
  D_FF_8 DFF_i_24 ( .D(s_D_Fmux_TFF[24]), .clk(clk), .Q(data_out[24]) );
  D_FF_7 DFF_i_25 ( .D(s_D_Fmux_TFF[25]), .clk(clk), .Q(data_out[25]) );
  D_FF_6 DFF_i_26 ( .D(s_D_Fmux_TFF[26]), .clk(clk), .Q(data_out[26]) );
  D_FF_5 DFF_i_27 ( .D(s_D_Fmux_TFF[27]), .clk(clk), .Q(data_out[27]) );
  D_FF_4 DFF_i_28 ( .D(s_D_Fmux_TFF[28]), .clk(clk), .Q(data_out[28]) );
  D_FF_3 DFF_i_29 ( .D(s_D_Fmux_TFF[29]), .clk(clk), .Q(data_out[29]) );
  D_FF_2 DFF_i_30 ( .D(s_D_Fmux_TFF[30]), .clk(clk), .Q(data_out[30]) );
  D_FF_1 DFF_i_31 ( .D(s_D_Fmux_TFF[31]), .clk(clk), .Q(data_out[31]) );
  Mux_Bit_NBIT_Sel2_0 MUX_0_0 ( .inputs({1'b0, data_out[0], data_out[31], 1'b0}), .sel({n7, n4}), .\output (s_D_Fmux_TFF[0]) );
  Mux_Bit_NBIT_Sel2_31 MUX_i_1 ( .inputs({1'b0, data_out[1:0], 1'b0}), .sel({
        n5, n2}), .\output (s_D_Fmux_TFF[1]) );
  Mux_Bit_NBIT_Sel2_30 MUX_i_2 ( .inputs({1'b0, data_out[2:1], 1'b0}), .sel({
        n5, n2}), .\output (s_D_Fmux_TFF[2]) );
  Mux_Bit_NBIT_Sel2_29 MUX_i_3 ( .inputs({1'b0, data_out[3:2], 1'b0}), .sel({
        n5, n2}), .\output (s_D_Fmux_TFF[3]) );
  Mux_Bit_NBIT_Sel2_28 MUX_i_4 ( .inputs({1'b0, data_out[4:3], 1'b0}), .sel({
        n5, n2}), .\output (s_D_Fmux_TFF[4]) );
  Mux_Bit_NBIT_Sel2_27 MUX_i_5 ( .inputs({1'b0, data_out[5:4], 1'b0}), .sel({
        n5, n2}), .\output (s_D_Fmux_TFF[5]) );
  Mux_Bit_NBIT_Sel2_26 MUX_i_6 ( .inputs({1'b0, data_out[6:5], 1'b0}), .sel({
        n5, n2}), .\output (s_D_Fmux_TFF[6]) );
  Mux_Bit_NBIT_Sel2_25 MUX_i_7 ( .inputs({1'b0, data_out[7:6], 1'b0}), .sel({
        n5, n2}), .\output (s_D_Fmux_TFF[7]) );
  Mux_Bit_NBIT_Sel2_24 MUX_i_8 ( .inputs({1'b0, data_out[8:7], 1'b0}), .sel({
        n5, n2}), .\output (s_D_Fmux_TFF[8]) );
  Mux_Bit_NBIT_Sel2_23 MUX_i_9 ( .inputs({1'b0, data_out[9:8], 1'b0}), .sel({
        n5, n2}), .\output (s_D_Fmux_TFF[9]) );
  Mux_Bit_NBIT_Sel2_22 MUX_i_10 ( .inputs({1'b0, data_out[10:9], 1'b0}), .sel(
        {n5, n2}), .\output (s_D_Fmux_TFF[10]) );
  Mux_Bit_NBIT_Sel2_21 MUX_i_11 ( .inputs({1'b0, data_out[11:10], 1'b0}), 
        .sel({n5, n2}), .\output (s_D_Fmux_TFF[11]) );
  Mux_Bit_NBIT_Sel2_20 MUX_i_12 ( .inputs({1'b0, data_out[12:11], 1'b0}), 
        .sel({n5, n2}), .\output (s_D_Fmux_TFF[12]) );
  Mux_Bit_NBIT_Sel2_19 MUX_i_13 ( .inputs({1'b0, data_out[13:12], 1'b0}), 
        .sel({n6, n3}), .\output (s_D_Fmux_TFF[13]) );
  Mux_Bit_NBIT_Sel2_18 MUX_i_14 ( .inputs({1'b0, data_out[14:13], 1'b0}), 
        .sel({n6, n3}), .\output (s_D_Fmux_TFF[14]) );
  Mux_Bit_NBIT_Sel2_17 MUX_i_15 ( .inputs({1'b0, data_out[15:14], 1'b0}), 
        .sel({n6, n3}), .\output (s_D_Fmux_TFF[15]) );
  Mux_Bit_NBIT_Sel2_16 MUX_i_16 ( .inputs({1'b0, data_out[16:15], 1'b0}), 
        .sel({n6, n3}), .\output (s_D_Fmux_TFF[16]) );
  Mux_Bit_NBIT_Sel2_15 MUX_i_17 ( .inputs({1'b0, data_out[17:16], 1'b0}), 
        .sel({n6, n3}), .\output (s_D_Fmux_TFF[17]) );
  Mux_Bit_NBIT_Sel2_14 MUX_i_18 ( .inputs({1'b0, data_out[18:17], 1'b0}), 
        .sel({n6, n3}), .\output (s_D_Fmux_TFF[18]) );
  Mux_Bit_NBIT_Sel2_13 MUX_i_19 ( .inputs({1'b0, data_out[19:18], 1'b0}), 
        .sel({n6, n3}), .\output (s_D_Fmux_TFF[19]) );
  Mux_Bit_NBIT_Sel2_12 MUX_i_20 ( .inputs({1'b0, data_out[20:19], 1'b0}), 
        .sel({n6, n3}), .\output (s_D_Fmux_TFF[20]) );
  Mux_Bit_NBIT_Sel2_11 MUX_i_21 ( .inputs({1'b0, data_out[21:20], 1'b0}), 
        .sel({n6, n3}), .\output (s_D_Fmux_TFF[21]) );
  Mux_Bit_NBIT_Sel2_10 MUX_i_22 ( .inputs({1'b0, data_out[22:21], 1'b0}), 
        .sel({n6, n3}), .\output (s_D_Fmux_TFF[22]) );
  Mux_Bit_NBIT_Sel2_9 MUX_i_23 ( .inputs({1'b0, data_out[23:22], 1'b0}), .sel(
        {n6, n3}), .\output (s_D_Fmux_TFF[23]) );
  Mux_Bit_NBIT_Sel2_8 MUX_i_24 ( .inputs({1'b0, data_out[24:23], 1'b0}), .sel(
        {n6, n3}), .\output (s_D_Fmux_TFF[24]) );
  Mux_Bit_NBIT_Sel2_7 MUX_i_25 ( .inputs({1'b0, data_out[25:24], 1'b0}), .sel(
        {n7, n4}), .\output (s_D_Fmux_TFF[25]) );
  Mux_Bit_NBIT_Sel2_6 MUX_i_26 ( .inputs({1'b0, data_out[26:25], 1'b0}), .sel(
        {n7, n4}), .\output (s_D_Fmux_TFF[26]) );
  Mux_Bit_NBIT_Sel2_5 MUX_i_27 ( .inputs({1'b0, data_out[27:26], 1'b0}), .sel(
        {n7, n4}), .\output (s_D_Fmux_TFF[27]) );
  Mux_Bit_NBIT_Sel2_4 MUX_i_28 ( .inputs({1'b0, data_out[28:27], 1'b0}), .sel(
        {n7, n4}), .\output (s_D_Fmux_TFF[28]) );
  Mux_Bit_NBIT_Sel2_3 MUX_i_29 ( .inputs({1'b0, data_out[29:28], 1'b0}), .sel(
        {n7, n4}), .\output (s_D_Fmux_TFF[29]) );
  Mux_Bit_NBIT_Sel2_2 MUX_i_30 ( .inputs({1'b0, data_out[30:29], 1'b0}), .sel(
        {n7, n4}), .\output (s_D_Fmux_TFF[30]) );
  Mux_Bit_NBIT_Sel2_1 MUX_i_31 ( .inputs({1'b1, data_out[31:30], 1'b1}), .sel(
        {n7, n4}), .\output (s_D_Fmux_TFF[31]) );
  BUF_X1 U3 ( .A(s_phi[0]), .Z(n4) );
  BUF_X1 U4 ( .A(s_phi[1]), .Z(n5) );
  BUF_X1 U5 ( .A(s_phi[1]), .Z(n6) );
  BUF_X1 U6 ( .A(s_phi[1]), .Z(n7) );
  BUF_X2 U7 ( .A(s_phi[0]), .Z(n2) );
  BUF_X2 U8 ( .A(s_phi[0]), .Z(n3) );
  AOI21_X1 U9 ( .B1(rotate), .B2(enable), .A(reset), .ZN(s_phi[1]) );
  AND3_X1 U10 ( .A1(rotate), .A2(n8), .A3(enable), .ZN(s_phi[0]) );
  INV_X1 U11 ( .A(reset), .ZN(n8) );
endmodule


module NPriorityEncoder_NBIT_OUT5 ( data_in, enable, data_out );
  input [31:0] data_in;
  output [4:0] data_out;
  input enable;
  wire   N369, N371, N373, N375, N377, n24, n25, n27, n28, n29, n30, n31, n32,
         n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46,
         n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60,
         n61, n62, n63, n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74,
         n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88,
         n89, n90, n91;

  DLH_X1 \data_out_reg[3]  ( .G(1'b1), .D(N375), .Q(data_out[3]) );
  DLH_X1 \data_out_reg[2]  ( .G(1'b1), .D(N373), .Q(data_out[2]) );
  DLH_X1 \data_out_reg[1]  ( .G(1'b1), .D(N371), .Q(data_out[1]) );
  DLH_X1 \data_out_reg[0]  ( .G(1'b1), .D(N369), .Q(data_out[0]) );
  NAND3_X1 U73 ( .A1(n51), .A2(n52), .A3(n53), .ZN(n50) );
  NAND3_X1 U74 ( .A1(n54), .A2(n55), .A3(n56), .ZN(n53) );
  NAND3_X1 U75 ( .A1(n62), .A2(n63), .A3(n64), .ZN(n61) );
  DLH_X1 \data_out_reg[4]  ( .G(1'b1), .D(N377), .Q(data_out[4]) );
  AOI21_X1 U3 ( .B1(n24), .B2(n25), .A(n91), .ZN(N377) );
  AND2_X1 U4 ( .A1(n31), .A2(n32), .ZN(n25) );
  NOR3_X1 U5 ( .A1(n48), .A2(data_in[25]), .A3(data_in[24]), .ZN(n45) );
  AOI211_X1 U6 ( .C1(n49), .C2(n50), .A(data_in[23]), .B(data_in[22]), .ZN(n48) );
  NOR2_X1 U8 ( .A1(data_in[21]), .A2(data_in[20]), .ZN(n49) );
  AOI21_X1 U9 ( .B1(n88), .B2(n62), .A(data_in[7]), .ZN(n86) );
  OAI21_X1 U10 ( .B1(data_in[4]), .B2(n89), .A(n66), .ZN(n88) );
  AOI21_X1 U11 ( .B1(data_in[1]), .B2(n90), .A(data_in[3]), .ZN(n89) );
  INV_X1 U12 ( .A(data_in[2]), .ZN(n90) );
  AOI21_X1 U13 ( .B1(n79), .B2(n51), .A(data_in[19]), .ZN(n77) );
  OAI21_X1 U14 ( .B1(data_in[16]), .B2(n80), .A(n55), .ZN(n79) );
  AOI21_X1 U15 ( .B1(n81), .B2(n58), .A(data_in[15]), .ZN(n80) );
  OAI21_X1 U16 ( .B1(data_in[12]), .B2(n82), .A(n83), .ZN(n81) );
  AOI21_X1 U17 ( .B1(n75), .B2(n76), .A(data_in[23]), .ZN(n73) );
  INV_X1 U18 ( .A(data_in[22]), .ZN(n76) );
  OAI21_X1 U19 ( .B1(data_in[20]), .B2(n77), .A(n78), .ZN(n75) );
  INV_X1 U20 ( .A(data_in[21]), .ZN(n78) );
  AOI21_X1 U21 ( .B1(n71), .B2(n72), .A(data_in[27]), .ZN(n70) );
  INV_X1 U22 ( .A(data_in[26]), .ZN(n72) );
  OAI21_X1 U23 ( .B1(data_in[24]), .B2(n73), .A(n74), .ZN(n71) );
  INV_X1 U24 ( .A(data_in[25]), .ZN(n74) );
  AOI21_X1 U25 ( .B1(n84), .B2(n85), .A(data_in[11]), .ZN(n82) );
  INV_X1 U26 ( .A(data_in[10]), .ZN(n85) );
  OAI21_X1 U27 ( .B1(data_in[8]), .B2(n86), .A(n87), .ZN(n84) );
  INV_X1 U28 ( .A(data_in[9]), .ZN(n87) );
  AOI21_X1 U29 ( .B1(n60), .B2(n61), .A(n30), .ZN(n57) );
  NOR2_X1 U30 ( .A1(data_in[9]), .A2(data_in[8]), .ZN(n60) );
  INV_X1 U31 ( .A(data_in[7]), .ZN(n63) );
  AOI21_X1 U32 ( .B1(n43), .B2(n44), .A(n91), .ZN(N371) );
  NOR2_X1 U33 ( .A1(data_in[31]), .A2(data_in[30]), .ZN(n43) );
  OAI211_X1 U34 ( .C1(n45), .C2(n46), .A(n34), .B(n47), .ZN(n44) );
  OR2_X1 U35 ( .A1(data_in[26]), .A2(data_in[27]), .ZN(n46) );
  OAI211_X1 U36 ( .C1(data_in[2]), .C2(data_in[3]), .A(n65), .B(n66), .ZN(n64)
         );
  INV_X1 U37 ( .A(data_in[4]), .ZN(n65) );
  OR2_X1 U38 ( .A1(data_in[11]), .A2(data_in[10]), .ZN(n30) );
  NOR2_X1 U39 ( .A1(n67), .A2(n91), .ZN(N369) );
  AOI21_X1 U40 ( .B1(n68), .B2(n69), .A(data_in[31]), .ZN(n67) );
  INV_X1 U41 ( .A(data_in[30]), .ZN(n69) );
  OAI21_X1 U42 ( .B1(data_in[28]), .B2(n70), .A(n47), .ZN(n68) );
  INV_X1 U43 ( .A(data_in[16]), .ZN(n54) );
  OAI211_X1 U44 ( .C1(n57), .C2(n41), .A(n58), .B(n59), .ZN(n56) );
  INV_X1 U45 ( .A(data_in[15]), .ZN(n59) );
  OR2_X1 U46 ( .A1(data_in[13]), .A2(data_in[12]), .ZN(n41) );
  INV_X1 U47 ( .A(data_in[14]), .ZN(n58) );
  INV_X1 U48 ( .A(data_in[5]), .ZN(n66) );
  INV_X1 U49 ( .A(data_in[18]), .ZN(n51) );
  INV_X1 U50 ( .A(data_in[6]), .ZN(n62) );
  INV_X1 U51 ( .A(data_in[17]), .ZN(n55) );
  INV_X1 U52 ( .A(data_in[13]), .ZN(n83) );
  INV_X1 U53 ( .A(data_in[19]), .ZN(n52) );
  NOR4_X1 U54 ( .A1(data_in[24]), .A2(data_in[25]), .A3(data_in[26]), .A4(
        data_in[27]), .ZN(n35) );
  NOR4_X1 U55 ( .A1(data_in[30]), .A2(data_in[31]), .A3(data_in[29]), .A4(n33), 
        .ZN(n24) );
  NAND2_X1 U56 ( .A1(n34), .A2(n35), .ZN(n33) );
  NOR4_X1 U57 ( .A1(data_in[16]), .A2(data_in[17]), .A3(data_in[18]), .A4(
        data_in[19]), .ZN(n32) );
  NOR4_X1 U58 ( .A1(data_in[20]), .A2(data_in[21]), .A3(data_in[22]), .A4(
        data_in[23]), .ZN(n31) );
  OAI21_X1 U59 ( .B1(n40), .B2(n29), .A(n32), .ZN(n39) );
  NOR4_X1 U60 ( .A1(data_in[9]), .A2(data_in[8]), .A3(n42), .A4(n30), .ZN(n40)
         );
  NOR4_X1 U61 ( .A1(data_in[7]), .A2(data_in[6]), .A3(data_in[5]), .A4(
        data_in[4]), .ZN(n42) );
  AOI21_X1 U62 ( .B1(n36), .B2(n37), .A(n91), .ZN(N373) );
  NOR3_X1 U63 ( .A1(data_in[29]), .A2(data_in[31]), .A3(data_in[30]), .ZN(n37)
         );
  AOI21_X1 U64 ( .B1(n35), .B2(n38), .A(data_in[28]), .ZN(n36) );
  NAND2_X1 U65 ( .A1(n31), .A2(n39), .ZN(n38) );
  AOI21_X1 U66 ( .B1(n24), .B2(n27), .A(n91), .ZN(N375) );
  NAND2_X1 U67 ( .A1(n25), .A2(n28), .ZN(n27) );
  OR4_X1 U68 ( .A1(n29), .A2(n30), .A3(data_in[8]), .A4(data_in[9]), .ZN(n28)
         );
  OR3_X1 U69 ( .A1(data_in[14]), .A2(data_in[15]), .A3(n41), .ZN(n29) );
  INV_X1 U70 ( .A(data_in[29]), .ZN(n47) );
  INV_X1 U71 ( .A(data_in[28]), .ZN(n34) );
  INV_X1 U72 ( .A(enable), .ZN(n91) );
endmodule


module ORGate_NX1_N32_0 ( A, B, Y );
  input [31:0] A;
  input [31:0] B;
  output Y;
  wire   n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20;

  NOR4_X1 U1 ( .A1(A[23]), .A2(A[22]), .A3(A[21]), .A4(A[20]), .ZN(n16) );
  NOR4_X1 U2 ( .A1(A[9]), .A2(A[8]), .A3(A[7]), .A4(A[6]), .ZN(n20) );
  NOR4_X1 U3 ( .A1(A[5]), .A2(A[4]), .A3(A[3]), .A4(A[31]), .ZN(n19) );
  NOR4_X1 U4 ( .A1(A[30]), .A2(A[2]), .A3(A[29]), .A4(A[28]), .ZN(n18) );
  NOR4_X1 U5 ( .A1(A[27]), .A2(A[26]), .A3(A[25]), .A4(A[24]), .ZN(n17) );
  NAND4_X1 U6 ( .A1(n13), .A2(n14), .A3(n15), .A4(n16), .ZN(n2) );
  NOR4_X1 U7 ( .A1(A[12]), .A2(A[11]), .A3(A[10]), .A4(A[0]), .ZN(n13) );
  NOR4_X1 U8 ( .A1(A[16]), .A2(A[15]), .A3(A[14]), .A4(A[13]), .ZN(n14) );
  NOR4_X1 U9 ( .A1(A[1]), .A2(A[19]), .A3(A[18]), .A4(A[17]), .ZN(n15) );
  OR4_X1 U10 ( .A1(n1), .A2(n2), .A3(n3), .A4(n4), .ZN(Y) );
  NAND4_X1 U11 ( .A1(n5), .A2(n6), .A3(n7), .A4(n8), .ZN(n4) );
  NAND4_X1 U12 ( .A1(n9), .A2(n10), .A3(n11), .A4(n12), .ZN(n3) );
  NAND4_X1 U13 ( .A1(n17), .A2(n18), .A3(n19), .A4(n20), .ZN(n1) );
  NOR4_X1 U14 ( .A1(B[9]), .A2(B[8]), .A3(B[7]), .A4(B[6]), .ZN(n12) );
  NOR4_X1 U15 ( .A1(B[23]), .A2(B[22]), .A3(B[21]), .A4(B[20]), .ZN(n8) );
  NOR4_X1 U16 ( .A1(B[5]), .A2(B[4]), .A3(B[3]), .A4(B[31]), .ZN(n11) );
  NOR4_X1 U17 ( .A1(B[1]), .A2(B[19]), .A3(B[18]), .A4(B[17]), .ZN(n7) );
  NOR4_X1 U18 ( .A1(B[30]), .A2(B[2]), .A3(B[29]), .A4(B[28]), .ZN(n10) );
  NOR4_X1 U19 ( .A1(B[16]), .A2(B[15]), .A3(B[14]), .A4(B[13]), .ZN(n6) );
  NOR4_X1 U20 ( .A1(B[27]), .A2(B[26]), .A3(B[25]), .A4(B[24]), .ZN(n9) );
  NOR4_X1 U21 ( .A1(B[12]), .A2(B[11]), .A3(B[10]), .A4(B[0]), .ZN(n5) );
endmodule


module NComparatorWithEnable_NBIT32_0 ( A, B, Enable, ComparatorBit );
  input [31:0] A;
  input [31:0] B;
  input Enable;
  output ComparatorBit;
  wire   \matrix[0][0] , \matrix[1][0] , \matrix[2][0] , \matrix[3][0] ,
         \matrix[4][0] , \matrix[5][0] , \matrix[6][0] , \matrix[7][0] ,
         \matrix[8][0] , \matrix[9][0] , \matrix[10][0] , \matrix[11][0] ,
         \matrix[12][0] , \matrix[13][0] , \matrix[14][0] , \matrix[15][0] ,
         \matrix[16][0] , \matrix[17][0] , \matrix[18][0] , \matrix[19][0] ,
         \matrix[20][0] , \matrix[21][0] , \matrix[22][0] , \matrix[23][0] ,
         \matrix[24][0] , \matrix[25][0] , \matrix[26][0] , \matrix[27][0] ,
         \matrix[28][0] , \matrix[29][0] , \matrix[30][0] , \matrix[31][0] ,
         n3, n1, n2, n4, n5, n6, n7, n8, n9, n10, n11, n14, n15, n16;
  assign n3 = Enable;

  ComparatorWithEnable_0 CWE_i_0 ( .a(A[0]), .b(B[0]), .enable(n16), .y(
        \matrix[0][0] ) );
  ComparatorWithEnable_1055 CWE_i_1 ( .a(A[1]), .b(B[1]), .enable(n14), .y(
        \matrix[1][0] ) );
  ComparatorWithEnable_1054 CWE_i_2 ( .a(A[2]), .b(B[2]), .enable(n14), .y(
        \matrix[2][0] ) );
  ComparatorWithEnable_1053 CWE_i_3 ( .a(A[3]), .b(B[3]), .enable(n14), .y(
        \matrix[3][0] ) );
  ComparatorWithEnable_1052 CWE_i_4 ( .a(A[4]), .b(B[4]), .enable(n14), .y(
        \matrix[4][0] ) );
  ComparatorWithEnable_1051 CWE_i_5 ( .a(A[5]), .b(B[5]), .enable(n14), .y(
        \matrix[5][0] ) );
  ComparatorWithEnable_1050 CWE_i_6 ( .a(A[6]), .b(B[6]), .enable(n14), .y(
        \matrix[6][0] ) );
  ComparatorWithEnable_1049 CWE_i_7 ( .a(A[7]), .b(B[7]), .enable(n14), .y(
        \matrix[7][0] ) );
  ComparatorWithEnable_1048 CWE_i_8 ( .a(A[8]), .b(B[8]), .enable(n14), .y(
        \matrix[8][0] ) );
  ComparatorWithEnable_1047 CWE_i_9 ( .a(A[9]), .b(B[9]), .enable(n14), .y(
        \matrix[9][0] ) );
  ComparatorWithEnable_1046 CWE_i_10 ( .a(A[10]), .b(B[10]), .enable(n14), .y(
        \matrix[10][0] ) );
  ComparatorWithEnable_1045 CWE_i_11 ( .a(A[11]), .b(B[11]), .enable(n14), .y(
        \matrix[11][0] ) );
  ComparatorWithEnable_1044 CWE_i_12 ( .a(A[12]), .b(B[12]), .enable(n14), .y(
        \matrix[12][0] ) );
  ComparatorWithEnable_1043 CWE_i_13 ( .a(A[13]), .b(B[13]), .enable(n15), .y(
        \matrix[13][0] ) );
  ComparatorWithEnable_1042 CWE_i_14 ( .a(A[14]), .b(B[14]), .enable(n15), .y(
        \matrix[14][0] ) );
  ComparatorWithEnable_1041 CWE_i_15 ( .a(A[15]), .b(B[15]), .enable(n15), .y(
        \matrix[15][0] ) );
  ComparatorWithEnable_1040 CWE_i_16 ( .a(A[16]), .b(B[16]), .enable(n15), .y(
        \matrix[16][0] ) );
  ComparatorWithEnable_1039 CWE_i_17 ( .a(A[17]), .b(B[17]), .enable(n15), .y(
        \matrix[17][0] ) );
  ComparatorWithEnable_1038 CWE_i_18 ( .a(A[18]), .b(B[18]), .enable(n15), .y(
        \matrix[18][0] ) );
  ComparatorWithEnable_1037 CWE_i_19 ( .a(A[19]), .b(B[19]), .enable(n15), .y(
        \matrix[19][0] ) );
  ComparatorWithEnable_1036 CWE_i_20 ( .a(A[20]), .b(B[20]), .enable(n15), .y(
        \matrix[20][0] ) );
  ComparatorWithEnable_1035 CWE_i_21 ( .a(A[21]), .b(B[21]), .enable(n15), .y(
        \matrix[21][0] ) );
  ComparatorWithEnable_1034 CWE_i_22 ( .a(A[22]), .b(B[22]), .enable(n15), .y(
        \matrix[22][0] ) );
  ComparatorWithEnable_1033 CWE_i_23 ( .a(A[23]), .b(B[23]), .enable(n15), .y(
        \matrix[23][0] ) );
  ComparatorWithEnable_1032 CWE_i_24 ( .a(A[24]), .b(B[24]), .enable(n15), .y(
        \matrix[24][0] ) );
  ComparatorWithEnable_1031 CWE_i_25 ( .a(A[25]), .b(B[25]), .enable(n16), .y(
        \matrix[25][0] ) );
  ComparatorWithEnable_1030 CWE_i_26 ( .a(A[26]), .b(B[26]), .enable(n16), .y(
        \matrix[26][0] ) );
  ComparatorWithEnable_1029 CWE_i_27 ( .a(A[27]), .b(B[27]), .enable(n16), .y(
        \matrix[27][0] ) );
  ComparatorWithEnable_1028 CWE_i_28 ( .a(A[28]), .b(B[28]), .enable(n16), .y(
        \matrix[28][0] ) );
  ComparatorWithEnable_1027 CWE_i_29 ( .a(A[29]), .b(B[29]), .enable(n16), .y(
        \matrix[29][0] ) );
  ComparatorWithEnable_1026 CWE_i_30 ( .a(A[30]), .b(B[30]), .enable(n16), .y(
        \matrix[30][0] ) );
  ComparatorWithEnable_1025 CWE_i_31 ( .a(A[31]), .b(B[31]), .enable(n16), .y(
        \matrix[31][0] ) );
  BUF_X1 U1 ( .A(n3), .Z(n15) );
  BUF_X1 U2 ( .A(n3), .Z(n14) );
  BUF_X1 U3 ( .A(n3), .Z(n16) );
  NAND4_X1 U4 ( .A1(\matrix[23][0] ), .A2(\matrix[22][0] ), .A3(
        \matrix[21][0] ), .A4(\matrix[20][0] ), .ZN(n7) );
  NAND4_X1 U5 ( .A1(\matrix[9][0] ), .A2(\matrix[8][0] ), .A3(\matrix[7][0] ), 
        .A4(\matrix[6][0] ), .ZN(n11) );
  NAND4_X1 U6 ( .A1(\matrix[1][0] ), .A2(\matrix[19][0] ), .A3(\matrix[18][0] ), .A4(\matrix[17][0] ), .ZN(n6) );
  NAND4_X1 U7 ( .A1(\matrix[5][0] ), .A2(\matrix[4][0] ), .A3(\matrix[3][0] ), 
        .A4(\matrix[31][0] ), .ZN(n10) );
  NAND4_X1 U8 ( .A1(\matrix[16][0] ), .A2(\matrix[15][0] ), .A3(
        \matrix[14][0] ), .A4(\matrix[13][0] ), .ZN(n5) );
  NAND4_X1 U9 ( .A1(\matrix[12][0] ), .A2(\matrix[11][0] ), .A3(
        \matrix[10][0] ), .A4(\matrix[0][0] ), .ZN(n4) );
  NAND4_X1 U10 ( .A1(\matrix[27][0] ), .A2(\matrix[26][0] ), .A3(
        \matrix[25][0] ), .A4(\matrix[24][0] ), .ZN(n8) );
  AND2_X1 U11 ( .A1(n1), .A2(n2), .ZN(ComparatorBit) );
  NOR4_X1 U12 ( .A1(n8), .A2(n9), .A3(n10), .A4(n11), .ZN(n1) );
  NOR4_X1 U13 ( .A1(n4), .A2(n5), .A3(n6), .A4(n7), .ZN(n2) );
  NAND4_X1 U14 ( .A1(\matrix[30][0] ), .A2(\matrix[2][0] ), .A3(
        \matrix[29][0] ), .A4(\matrix[28][0] ), .ZN(n9) );
endmodule


module Mux_1Bit_2X1_6 ( port0, port1, sel, portY );
  input port0, port1, sel;
  output portY;
  wire   n3, n4;

  INV_X1 U1 ( .A(n3), .ZN(portY) );
  AOI22_X1 U2 ( .A1(port0), .A2(n4), .B1(sel), .B2(port1), .ZN(n3) );
  INV_X1 U3 ( .A(sel), .ZN(n4) );
endmodule


module Mux_1Bit_2X1_0 ( port0, port1, sel, portY );
  input port0, port1, sel;
  output portY;
  wire   n3, n1;

  INV_X1 U1 ( .A(n3), .ZN(portY) );
  AOI22_X1 U2 ( .A1(port0), .A2(n1), .B1(sel), .B2(port1), .ZN(n3) );
  INV_X1 U3 ( .A(sel), .ZN(n1) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_127 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  INV_X1 U1 ( .A(n14), .ZN(n4) );
  INV_X1 U2 ( .A(n14), .ZN(n5) );
  BUF_X1 U3 ( .A(n2), .Z(n11) );
  BUF_X1 U4 ( .A(n3), .Z(n12) );
  BUF_X1 U5 ( .A(n1), .Z(n6) );
  BUF_X1 U6 ( .A(n2), .Z(n10) );
  BUF_X1 U7 ( .A(n1), .Z(n7) );
  BUF_X1 U8 ( .A(n2), .Z(n9) );
  BUF_X1 U9 ( .A(n1), .Z(n8) );
  BUF_X1 U10 ( .A(n3), .Z(n14) );
  BUF_X1 U11 ( .A(n3), .Z(n13) );
  BUF_X1 U12 ( .A(sel), .Z(n3) );
  BUF_X1 U13 ( .A(sel), .Z(n2) );
  BUF_X1 U14 ( .A(sel), .Z(n1) );
  INV_X1 U15 ( .A(n53), .ZN(N22) );
  AOI22_X1 U16 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n10), .ZN(n53)
         );
  INV_X1 U17 ( .A(n52), .ZN(N23) );
  AOI22_X1 U18 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n9), .ZN(n52) );
  INV_X1 U19 ( .A(n51), .ZN(N24) );
  AOI22_X1 U20 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n9), .ZN(n51) );
  INV_X1 U21 ( .A(n50), .ZN(N25) );
  AOI22_X1 U22 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n9), .ZN(n50) );
  INV_X1 U23 ( .A(n57), .ZN(N19) );
  AOI22_X1 U24 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n11), .ZN(n57)
         );
  INV_X1 U25 ( .A(n55), .ZN(N20) );
  AOI22_X1 U26 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n10), .ZN(n55)
         );
  INV_X1 U27 ( .A(n54), .ZN(N21) );
  AOI22_X1 U28 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n10), .ZN(n54)
         );
  INV_X1 U29 ( .A(n45), .ZN(N3) );
  AOI22_X1 U30 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n8), .ZN(n45) );
  INV_X1 U31 ( .A(n61), .ZN(N15) );
  AOI22_X1 U32 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n12), .ZN(n61)
         );
  INV_X1 U33 ( .A(n60), .ZN(N16) );
  AOI22_X1 U34 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n12), .ZN(n60)
         );
  INV_X1 U35 ( .A(n59), .ZN(N17) );
  AOI22_X1 U36 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n11), .ZN(n59)
         );
  INV_X1 U37 ( .A(n58), .ZN(N18) );
  AOI22_X1 U38 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n11), .ZN(n58)
         );
  INV_X1 U39 ( .A(n56), .ZN(N2) );
  AOI22_X1 U40 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n11), .ZN(n56) );
  INV_X1 U41 ( .A(n64), .ZN(N12) );
  AOI22_X1 U42 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n13), .ZN(n64)
         );
  INV_X1 U43 ( .A(n63), .ZN(N13) );
  AOI22_X1 U44 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n12), .ZN(n63)
         );
  INV_X1 U45 ( .A(n62), .ZN(N14) );
  AOI22_X1 U46 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n12), .ZN(n62)
         );
  INV_X1 U47 ( .A(n36), .ZN(N8) );
  AOI22_X1 U48 ( .A1(port0[6]), .A2(n4), .B1(port1[6]), .B2(n6), .ZN(n36) );
  INV_X1 U49 ( .A(n34), .ZN(N9) );
  AOI22_X1 U50 ( .A1(port0[7]), .A2(n5), .B1(n13), .B2(port1[7]), .ZN(n34) );
  INV_X1 U51 ( .A(n66), .ZN(N10) );
  AOI22_X1 U52 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n13), .ZN(n66) );
  INV_X1 U53 ( .A(n65), .ZN(N11) );
  AOI22_X1 U54 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n13), .ZN(n65) );
  INV_X1 U55 ( .A(n39), .ZN(N5) );
  AOI22_X1 U56 ( .A1(port0[3]), .A2(n5), .B1(port1[3]), .B2(n6), .ZN(n39) );
  INV_X1 U57 ( .A(n38), .ZN(N6) );
  AOI22_X1 U58 ( .A1(port0[4]), .A2(n4), .B1(port1[4]), .B2(n6), .ZN(n38) );
  INV_X1 U59 ( .A(n41), .ZN(N33) );
  AOI22_X1 U60 ( .A1(port0[31]), .A2(n4), .B1(port1[31]), .B2(n7), .ZN(n41) );
  INV_X1 U61 ( .A(n37), .ZN(N7) );
  AOI22_X1 U62 ( .A1(port0[5]), .A2(n5), .B1(port1[5]), .B2(n6), .ZN(n37) );
  INV_X1 U63 ( .A(n40), .ZN(N4) );
  AOI22_X1 U64 ( .A1(port0[2]), .A2(n4), .B1(port1[2]), .B2(n7), .ZN(n40) );
  INV_X1 U65 ( .A(n44), .ZN(N30) );
  AOI22_X1 U66 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n7), .ZN(n44) );
  INV_X1 U67 ( .A(n43), .ZN(N31) );
  AOI22_X1 U68 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n10), .ZN(n43)
         );
  INV_X1 U69 ( .A(n42), .ZN(N32) );
  AOI22_X1 U70 ( .A1(port0[30]), .A2(n5), .B1(port1[30]), .B2(n7), .ZN(n42) );
  INV_X1 U71 ( .A(n49), .ZN(N26) );
  AOI22_X1 U72 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n9), .ZN(n49) );
  INV_X1 U73 ( .A(n48), .ZN(N27) );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n8), .ZN(n48) );
  INV_X1 U75 ( .A(n47), .ZN(N28) );
  AOI22_X1 U76 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n8), .ZN(n47) );
  INV_X1 U77 ( .A(n46), .ZN(N29) );
  AOI22_X1 U78 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n8), .ZN(n46) );
endmodule


module SAT_Counter_N2 ( SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, 
        SAT_setToDef, SAT_SO );
  output [1:0] SAT_SO;
  input SAT_clk, SAT_reset, SAT_enable, SAT_Ud, SAT_update, SAT_setToDef;
  wire   s_enable, s_Ud, s_clk, s_reset, s_TcMax, s_TcMin;

  UD_COUNTER_UDC_NBIT2 CNT ( .UDC_EN(s_enable), .UDC_UP(s_Ud), .UDC_CLK(s_clk), 
        .UDC_RST(s_reset), .UDC_OUT(SAT_SO) );
  CU_SatCounter_0 CU ( .CU_clk(SAT_clk), .CU_reset(SAT_reset), .CU_enable(
        SAT_enable), .CU_Ud(SAT_Ud), .CU_update(SAT_update), .CU_loadDefault(
        SAT_setToDef), .CU_TcMax(s_TcMax), .CU_TcMin(s_TcMin), .UDC_clk(s_clk), 
        .UDC_Ud(s_Ud), .UDC_enable(s_enable), .UDC_reset(s_reset) );
  ANDGate_NX1_N2 AND1 ( .A(SAT_SO), .B({1'b1, 1'b1}), .Y(s_TcMax) );
  NORGate_NX1_N2 NOR1 ( .A(SAT_SO), .B({1'b0, 1'b0}), .Y(s_TcMin) );
endmodule


module NRegister_N4 ( clk, reset, data_in, enable, load, data_out );
  input [3:0] data_in;
  output [3:0] data_out;
  input clk, reset, enable, load;
  wire   n12, n13, n14, n16, n1, n2, n3, net106788, n10, n11, n17, n18, n19,
         n20, n5;

  DFFR_X1 \data_out_reg[0]  ( .D(n12), .CK(clk), .RN(n5), .Q(data_out[0]), 
        .QN(net106788) );
  DFFR_X1 \data_out_reg[3]  ( .D(n16), .CK(clk), .RN(n5), .Q(data_out[3]), 
        .QN(n2) );
  DFFR_X1 \data_out_reg[2]  ( .D(n14), .CK(clk), .RN(n5), .Q(data_out[2]), 
        .QN(n1) );
  DFFR_X1 \data_out_reg[1]  ( .D(n13), .CK(clk), .RN(n5), .Q(data_out[1]), 
        .QN(n3) );
  INV_X1 U3 ( .A(n10), .ZN(n17) );
  NAND2_X1 U4 ( .A1(load), .A2(enable), .ZN(n10) );
  OAI22_X1 U5 ( .A1(n10), .A2(n18), .B1(n1), .B2(n17), .ZN(n14) );
  INV_X1 U6 ( .A(data_in[2]), .ZN(n18) );
  OAI22_X1 U7 ( .A1(n10), .A2(n19), .B1(n3), .B2(n17), .ZN(n13) );
  INV_X1 U8 ( .A(data_in[1]), .ZN(n19) );
  OAI22_X1 U9 ( .A1(n10), .A2(n11), .B1(n2), .B2(n17), .ZN(n16) );
  INV_X1 U10 ( .A(data_in[3]), .ZN(n11) );
  OAI22_X1 U11 ( .A1(n10), .A2(n20), .B1(net106788), .B2(n17), .ZN(n12) );
  INV_X1 U12 ( .A(data_in[0]), .ZN(n20) );
  INV_X1 U13 ( .A(reset), .ZN(n5) );
endmodule


module NRegister_N10 ( clk, reset, data_in, enable, load, data_out );
  input [9:0] data_in;
  output [9:0] data_out;
  input clk, reset, enable, load;
  wire   n24, n25, n26, n27, n28, n29, n30, n31, n32, n34, n1, n2, n3,
         net106782, net106783, net106784, net106785, net106786, net106787, n17,
         n18, n19, n20, n21, n22, n23, n35, n36, n37, n38, n39, n8;

  DFFR_X1 \data_out_reg[8]  ( .D(n32), .CK(clk), .RN(n8), .Q(data_out[8]) );
  DFFR_X1 \data_out_reg[7]  ( .D(n31), .CK(clk), .RN(n8), .Q(data_out[7]), 
        .QN(net106787) );
  DFFR_X1 \data_out_reg[6]  ( .D(n30), .CK(clk), .RN(n8), .Q(data_out[6]), 
        .QN(net106786) );
  DFFR_X1 \data_out_reg[3]  ( .D(n27), .CK(clk), .RN(n8), .Q(data_out[3]), 
        .QN(net106785) );
  DFFR_X1 \data_out_reg[2]  ( .D(n26), .CK(clk), .RN(n8), .Q(data_out[2]), 
        .QN(net106784) );
  DFFR_X1 \data_out_reg[1]  ( .D(n25), .CK(clk), .RN(n8), .Q(data_out[1]), 
        .QN(net106783) );
  DFFR_X1 \data_out_reg[0]  ( .D(n24), .CK(clk), .RN(n8), .Q(data_out[0]), 
        .QN(net106782) );
  DFFR_X1 \data_out_reg[4]  ( .D(n28), .CK(clk), .RN(n8), .Q(data_out[4]), 
        .QN(n2) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n8), .Q(data_out[5]), 
        .QN(n1) );
  DFFR_X1 \data_out_reg[9]  ( .D(n34), .CK(clk), .RN(n8), .Q(data_out[9]), 
        .QN(n3) );
  INV_X1 U3 ( .A(n17), .ZN(n19) );
  NAND2_X1 U4 ( .A1(load), .A2(enable), .ZN(n17) );
  OAI22_X1 U5 ( .A1(n17), .A2(n23), .B1(n1), .B2(n19), .ZN(n29) );
  INV_X1 U6 ( .A(data_in[5]), .ZN(n23) );
  OAI22_X1 U7 ( .A1(n17), .A2(n35), .B1(n2), .B2(n19), .ZN(n28) );
  INV_X1 U8 ( .A(data_in[4]), .ZN(n35) );
  OAI22_X1 U9 ( .A1(n17), .A2(n18), .B1(n3), .B2(n19), .ZN(n34) );
  INV_X1 U10 ( .A(data_in[9]), .ZN(n18) );
  OAI22_X1 U11 ( .A1(n17), .A2(n39), .B1(net106782), .B2(n19), .ZN(n24) );
  INV_X1 U12 ( .A(data_in[0]), .ZN(n39) );
  OAI22_X1 U13 ( .A1(n17), .A2(n38), .B1(net106783), .B2(n19), .ZN(n25) );
  INV_X1 U14 ( .A(data_in[1]), .ZN(n38) );
  OAI22_X1 U15 ( .A1(n17), .A2(n37), .B1(net106784), .B2(n19), .ZN(n26) );
  INV_X1 U16 ( .A(data_in[2]), .ZN(n37) );
  OAI22_X1 U17 ( .A1(n17), .A2(n36), .B1(net106785), .B2(n19), .ZN(n27) );
  INV_X1 U18 ( .A(data_in[3]), .ZN(n36) );
  OAI22_X1 U19 ( .A1(n17), .A2(n22), .B1(net106786), .B2(n19), .ZN(n30) );
  INV_X1 U20 ( .A(data_in[6]), .ZN(n22) );
  OAI22_X1 U21 ( .A1(n17), .A2(n21), .B1(net106787), .B2(n19), .ZN(n31) );
  INV_X1 U22 ( .A(data_in[7]), .ZN(n21) );
  INV_X1 U23 ( .A(n20), .ZN(n32) );
  AOI22_X1 U24 ( .A1(n19), .A2(data_in[8]), .B1(n17), .B2(data_out[8]), .ZN(
        n20) );
  INV_X1 U25 ( .A(reset), .ZN(n8) );
endmodule


module NRegister_N19 ( clk, reset, data_in, enable, load, data_out );
  input [18:0] data_in;
  output [18:0] data_out;
  input clk, reset, enable, load;
  wire   n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n61, n1, net106767, net106768, net106769,
         net106770, net106771, net106772, net106773, net106774, net106775,
         net106776, net106777, net106778, net106779, net106780, net106781, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n62, n63, n64,
         n65, n66, n67, n68, n69, n70, n12, n13;

  DFFR_X1 \data_out_reg[18]  ( .D(n61), .CK(clk), .RN(n13), .Q(data_out[18]), 
        .QN(net106781) );
  DFFR_X1 \data_out_reg[17]  ( .D(n59), .CK(clk), .RN(n13), .Q(data_out[17])
         );
  DFFR_X1 \data_out_reg[15]  ( .D(n57), .CK(clk), .RN(n13), .Q(data_out[15])
         );
  DFFR_X1 \data_out_reg[14]  ( .D(n56), .CK(clk), .RN(n13), .Q(data_out[14]), 
        .QN(net106780) );
  DFFR_X1 \data_out_reg[13]  ( .D(n55), .CK(clk), .RN(n13), .Q(data_out[13]), 
        .QN(net106779) );
  DFFR_X1 \data_out_reg[12]  ( .D(n54), .CK(clk), .RN(n13), .Q(data_out[12])
         );
  DFFR_X1 \data_out_reg[11]  ( .D(n53), .CK(clk), .RN(n13), .Q(data_out[11]), 
        .QN(net106778) );
  DFFR_X1 \data_out_reg[10]  ( .D(n52), .CK(clk), .RN(n13), .Q(data_out[10]), 
        .QN(net106777) );
  DFFR_X1 \data_out_reg[9]  ( .D(n51), .CK(clk), .RN(n13), .Q(data_out[9]), 
        .QN(net106776) );
  DFFR_X1 \data_out_reg[8]  ( .D(n50), .CK(clk), .RN(n13), .Q(data_out[8]), 
        .QN(net106775) );
  DFFR_X1 \data_out_reg[7]  ( .D(n49), .CK(clk), .RN(n13), .Q(data_out[7]), 
        .QN(net106774) );
  DFFR_X1 \data_out_reg[6]  ( .D(n48), .CK(clk), .RN(n13), .Q(data_out[6]), 
        .QN(net106773) );
  DFFR_X1 \data_out_reg[5]  ( .D(n47), .CK(clk), .RN(n13), .Q(data_out[5]), 
        .QN(net106772) );
  DFFR_X1 \data_out_reg[4]  ( .D(n46), .CK(clk), .RN(n13), .Q(data_out[4]), 
        .QN(net106771) );
  DFFR_X1 \data_out_reg[3]  ( .D(n45), .CK(clk), .RN(n13), .Q(data_out[3]), 
        .QN(net106770) );
  DFFR_X1 \data_out_reg[2]  ( .D(n44), .CK(clk), .RN(n13), .Q(data_out[2]), 
        .QN(net106769) );
  DFFR_X1 \data_out_reg[1]  ( .D(n43), .CK(clk), .RN(n13), .Q(data_out[1]), 
        .QN(net106768) );
  DFFR_X1 \data_out_reg[0]  ( .D(n42), .CK(clk), .RN(n13), .Q(data_out[0]), 
        .QN(net106767) );
  DFFR_X1 \data_out_reg[16]  ( .D(n58), .CK(clk), .RN(n13), .Q(data_out[16]), 
        .QN(n1) );
  INV_X1 U3 ( .A(n30), .ZN(n32) );
  NAND2_X1 U4 ( .A1(load), .A2(enable), .ZN(n30) );
  NAND2_X1 U5 ( .A1(load), .A2(enable), .ZN(n12) );
  OAI22_X1 U6 ( .A1(n30), .A2(n34), .B1(n1), .B2(n32), .ZN(n58) );
  INV_X1 U7 ( .A(data_in[16]), .ZN(n34) );
  OAI22_X1 U8 ( .A1(n30), .A2(n70), .B1(net106767), .B2(n32), .ZN(n42) );
  INV_X1 U9 ( .A(data_in[0]), .ZN(n70) );
  OAI22_X1 U10 ( .A1(n12), .A2(n69), .B1(net106768), .B2(n32), .ZN(n43) );
  INV_X1 U11 ( .A(data_in[1]), .ZN(n69) );
  OAI22_X1 U12 ( .A1(n30), .A2(n68), .B1(net106769), .B2(n32), .ZN(n44) );
  INV_X1 U13 ( .A(data_in[2]), .ZN(n68) );
  OAI22_X1 U14 ( .A1(n12), .A2(n67), .B1(net106770), .B2(n32), .ZN(n45) );
  INV_X1 U15 ( .A(data_in[3]), .ZN(n67) );
  OAI22_X1 U16 ( .A1(n30), .A2(n66), .B1(net106771), .B2(n32), .ZN(n46) );
  INV_X1 U17 ( .A(data_in[4]), .ZN(n66) );
  OAI22_X1 U18 ( .A1(n12), .A2(n65), .B1(net106772), .B2(n32), .ZN(n47) );
  INV_X1 U19 ( .A(data_in[5]), .ZN(n65) );
  OAI22_X1 U20 ( .A1(n30), .A2(n64), .B1(net106773), .B2(n32), .ZN(n48) );
  INV_X1 U21 ( .A(data_in[6]), .ZN(n64) );
  OAI22_X1 U22 ( .A1(n12), .A2(n63), .B1(net106774), .B2(n32), .ZN(n49) );
  INV_X1 U23 ( .A(data_in[7]), .ZN(n63) );
  OAI22_X1 U24 ( .A1(n30), .A2(n62), .B1(net106775), .B2(n32), .ZN(n50) );
  INV_X1 U25 ( .A(data_in[8]), .ZN(n62) );
  OAI22_X1 U26 ( .A1(n12), .A2(n41), .B1(net106776), .B2(n32), .ZN(n51) );
  INV_X1 U27 ( .A(data_in[9]), .ZN(n41) );
  OAI22_X1 U28 ( .A1(n30), .A2(n40), .B1(net106777), .B2(n32), .ZN(n52) );
  INV_X1 U29 ( .A(data_in[10]), .ZN(n40) );
  OAI22_X1 U30 ( .A1(n12), .A2(n39), .B1(net106778), .B2(n32), .ZN(n53) );
  INV_X1 U31 ( .A(data_in[11]), .ZN(n39) );
  OAI22_X1 U32 ( .A1(n30), .A2(n37), .B1(net106779), .B2(n32), .ZN(n55) );
  INV_X1 U33 ( .A(data_in[13]), .ZN(n37) );
  OAI22_X1 U34 ( .A1(n12), .A2(n36), .B1(net106780), .B2(n32), .ZN(n56) );
  INV_X1 U35 ( .A(data_in[14]), .ZN(n36) );
  OAI22_X1 U36 ( .A1(n12), .A2(n31), .B1(net106781), .B2(n32), .ZN(n61) );
  INV_X1 U37 ( .A(data_in[18]), .ZN(n31) );
  INV_X1 U38 ( .A(n38), .ZN(n54) );
  AOI22_X1 U39 ( .A1(n32), .A2(data_in[12]), .B1(data_out[12]), .B2(n12), .ZN(
        n38) );
  INV_X1 U40 ( .A(n35), .ZN(n57) );
  AOI22_X1 U41 ( .A1(n32), .A2(data_in[15]), .B1(data_out[15]), .B2(n30), .ZN(
        n35) );
  INV_X1 U42 ( .A(n33), .ZN(n59) );
  AOI22_X1 U43 ( .A1(n32), .A2(data_in[17]), .B1(n12), .B2(data_out[17]), .ZN(
        n33) );
  INV_X1 U44 ( .A(reset), .ZN(n13) );
endmodule


module NRegister_N26 ( clk, reset, data_in, enable, load, data_out );
  input [25:0] data_in;
  output [25:0] data_out;
  input clk, reset, enable, load;
  wire   n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n82, net106741,
         net106742, net106743, net106744, net106745, net106746, net106747,
         net106748, net106749, net106750, net106751, net106752, net106753,
         net106754, net106755, net106756, net106757, net106758, net106759,
         net106760, net106761, net106762, net106763, net106764, net106765,
         net106766, n29, n30, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41,
         n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54, n55,
         n83, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  DFFR_X1 \data_out_reg[25]  ( .D(n82), .CK(clk), .RN(n12), .Q(data_out[25]), 
        .QN(net106766) );
  DFFR_X1 \data_out_reg[24]  ( .D(n80), .CK(clk), .RN(n12), .Q(data_out[24]), 
        .QN(net106765) );
  DFFR_X1 \data_out_reg[23]  ( .D(n79), .CK(clk), .RN(n12), .Q(data_out[23]), 
        .QN(net106764) );
  DFFR_X1 \data_out_reg[22]  ( .D(n78), .CK(clk), .RN(n12), .Q(data_out[22]), 
        .QN(net106763) );
  DFFR_X1 \data_out_reg[21]  ( .D(n77), .CK(clk), .RN(n12), .Q(data_out[21]), 
        .QN(net106762) );
  DFFR_X1 \data_out_reg[20]  ( .D(n76), .CK(clk), .RN(n12), .Q(data_out[20]), 
        .QN(net106761) );
  DFFR_X1 \data_out_reg[19]  ( .D(n75), .CK(clk), .RN(n13), .Q(data_out[19]), 
        .QN(net106760) );
  DFFR_X1 \data_out_reg[18]  ( .D(n74), .CK(clk), .RN(n11), .Q(data_out[18]), 
        .QN(net106759) );
  DFFR_X1 \data_out_reg[17]  ( .D(n73), .CK(clk), .RN(n11), .Q(data_out[17]), 
        .QN(net106758) );
  DFFR_X1 \data_out_reg[16]  ( .D(n72), .CK(clk), .RN(n11), .Q(data_out[16]), 
        .QN(net106757) );
  DFFR_X1 \data_out_reg[15]  ( .D(n71), .CK(clk), .RN(n11), .Q(data_out[15]), 
        .QN(net106756) );
  DFFR_X1 \data_out_reg[14]  ( .D(n70), .CK(clk), .RN(n11), .Q(data_out[14]), 
        .QN(net106755) );
  DFFR_X1 \data_out_reg[13]  ( .D(n69), .CK(clk), .RN(n11), .Q(data_out[13]), 
        .QN(net106754) );
  DFFR_X1 \data_out_reg[12]  ( .D(n68), .CK(clk), .RN(n11), .Q(data_out[12]), 
        .QN(net106753) );
  DFFR_X1 \data_out_reg[11]  ( .D(n67), .CK(clk), .RN(n11), .Q(data_out[11]), 
        .QN(net106752) );
  DFFR_X1 \data_out_reg[10]  ( .D(n66), .CK(clk), .RN(n11), .Q(data_out[10]), 
        .QN(net106751) );
  DFFR_X1 \data_out_reg[9]  ( .D(n65), .CK(clk), .RN(n11), .Q(data_out[9]), 
        .QN(net106750) );
  DFFR_X1 \data_out_reg[8]  ( .D(n64), .CK(clk), .RN(n11), .Q(data_out[8]), 
        .QN(net106749) );
  DFFR_X1 \data_out_reg[7]  ( .D(n63), .CK(clk), .RN(n13), .Q(data_out[7]), 
        .QN(net106748) );
  DFFR_X1 \data_out_reg[6]  ( .D(n62), .CK(clk), .RN(n12), .Q(data_out[6]), 
        .QN(net106747) );
  DFFR_X1 \data_out_reg[5]  ( .D(n61), .CK(clk), .RN(n12), .Q(data_out[5]), 
        .QN(net106746) );
  DFFR_X1 \data_out_reg[4]  ( .D(n60), .CK(clk), .RN(n12), .Q(data_out[4]), 
        .QN(net106745) );
  DFFR_X1 \data_out_reg[3]  ( .D(n59), .CK(clk), .RN(n12), .Q(data_out[3]), 
        .QN(net106744) );
  DFFR_X1 \data_out_reg[2]  ( .D(n58), .CK(clk), .RN(n12), .Q(data_out[2]), 
        .QN(net106743) );
  DFFR_X1 \data_out_reg[1]  ( .D(n57), .CK(clk), .RN(n12), .Q(data_out[1]), 
        .QN(net106742) );
  DFFR_X1 \data_out_reg[0]  ( .D(n56), .CK(clk), .RN(n11), .Q(data_out[0]), 
        .QN(net106741) );
  INV_X1 U3 ( .A(n7), .ZN(n10) );
  BUF_X1 U4 ( .A(n8), .Z(n6) );
  BUF_X1 U5 ( .A(n8), .Z(n5) );
  BUF_X1 U6 ( .A(n9), .Z(n4) );
  BUF_X1 U7 ( .A(n9), .Z(n3) );
  BUF_X1 U8 ( .A(n9), .Z(n2) );
  BUF_X1 U9 ( .A(n8), .Z(n7) );
  BUF_X1 U10 ( .A(n29), .Z(n8) );
  BUF_X1 U11 ( .A(n29), .Z(n9) );
  BUF_X1 U12 ( .A(n14), .Z(n11) );
  BUF_X1 U13 ( .A(n14), .Z(n12) );
  BUF_X1 U14 ( .A(n14), .Z(n13) );
  OAI22_X1 U15 ( .A1(n7), .A2(n83), .B1(net106741), .B2(n10), .ZN(n56) );
  INV_X1 U16 ( .A(data_in[0]), .ZN(n83) );
  OAI22_X1 U17 ( .A1(n6), .A2(n55), .B1(net106742), .B2(n10), .ZN(n57) );
  INV_X1 U18 ( .A(data_in[1]), .ZN(n55) );
  OAI22_X1 U19 ( .A1(n6), .A2(n54), .B1(net106743), .B2(n10), .ZN(n58) );
  INV_X1 U20 ( .A(data_in[2]), .ZN(n54) );
  OAI22_X1 U21 ( .A1(n6), .A2(n53), .B1(net106744), .B2(n10), .ZN(n59) );
  INV_X1 U22 ( .A(data_in[3]), .ZN(n53) );
  OAI22_X1 U23 ( .A1(n6), .A2(n52), .B1(net106745), .B2(n10), .ZN(n60) );
  INV_X1 U24 ( .A(data_in[4]), .ZN(n52) );
  OAI22_X1 U25 ( .A1(n6), .A2(n51), .B1(net106746), .B2(n10), .ZN(n61) );
  INV_X1 U26 ( .A(data_in[5]), .ZN(n51) );
  OAI22_X1 U27 ( .A1(n5), .A2(n50), .B1(net106747), .B2(n10), .ZN(n62) );
  INV_X1 U28 ( .A(data_in[6]), .ZN(n50) );
  OAI22_X1 U29 ( .A1(n5), .A2(n49), .B1(net106748), .B2(n10), .ZN(n63) );
  INV_X1 U30 ( .A(data_in[7]), .ZN(n49) );
  OAI22_X1 U31 ( .A1(n5), .A2(n48), .B1(net106749), .B2(n10), .ZN(n64) );
  INV_X1 U32 ( .A(data_in[8]), .ZN(n48) );
  OAI22_X1 U33 ( .A1(n5), .A2(n47), .B1(net106750), .B2(n10), .ZN(n65) );
  INV_X1 U34 ( .A(data_in[9]), .ZN(n47) );
  OAI22_X1 U35 ( .A1(n5), .A2(n46), .B1(net106751), .B2(n10), .ZN(n66) );
  INV_X1 U36 ( .A(data_in[10]), .ZN(n46) );
  OAI22_X1 U37 ( .A1(n4), .A2(n45), .B1(net106752), .B2(n10), .ZN(n67) );
  INV_X1 U38 ( .A(data_in[11]), .ZN(n45) );
  OAI22_X1 U39 ( .A1(n4), .A2(n44), .B1(net106753), .B2(n10), .ZN(n68) );
  INV_X1 U40 ( .A(data_in[12]), .ZN(n44) );
  OAI22_X1 U41 ( .A1(n4), .A2(n43), .B1(net106754), .B2(n10), .ZN(n69) );
  INV_X1 U42 ( .A(data_in[13]), .ZN(n43) );
  OAI22_X1 U43 ( .A1(n4), .A2(n42), .B1(net106755), .B2(n10), .ZN(n70) );
  INV_X1 U44 ( .A(data_in[14]), .ZN(n42) );
  OAI22_X1 U45 ( .A1(n4), .A2(n41), .B1(net106756), .B2(n10), .ZN(n71) );
  INV_X1 U46 ( .A(data_in[15]), .ZN(n41) );
  OAI22_X1 U47 ( .A1(n3), .A2(n40), .B1(net106757), .B2(n10), .ZN(n72) );
  INV_X1 U48 ( .A(data_in[16]), .ZN(n40) );
  OAI22_X1 U49 ( .A1(n3), .A2(n39), .B1(net106758), .B2(n10), .ZN(n73) );
  INV_X1 U50 ( .A(data_in[17]), .ZN(n39) );
  OAI22_X1 U51 ( .A1(n3), .A2(n38), .B1(net106759), .B2(n10), .ZN(n74) );
  INV_X1 U52 ( .A(data_in[18]), .ZN(n38) );
  OAI22_X1 U53 ( .A1(n3), .A2(n37), .B1(net106760), .B2(n10), .ZN(n75) );
  INV_X1 U54 ( .A(data_in[19]), .ZN(n37) );
  OAI22_X1 U55 ( .A1(n3), .A2(n36), .B1(net106761), .B2(n10), .ZN(n76) );
  INV_X1 U56 ( .A(data_in[20]), .ZN(n36) );
  OAI22_X1 U57 ( .A1(n2), .A2(n35), .B1(net106762), .B2(n10), .ZN(n77) );
  INV_X1 U58 ( .A(data_in[21]), .ZN(n35) );
  OAI22_X1 U59 ( .A1(n2), .A2(n34), .B1(net106763), .B2(n10), .ZN(n78) );
  INV_X1 U60 ( .A(data_in[22]), .ZN(n34) );
  OAI22_X1 U61 ( .A1(n2), .A2(n33), .B1(net106764), .B2(n10), .ZN(n79) );
  INV_X1 U62 ( .A(data_in[23]), .ZN(n33) );
  OAI22_X1 U63 ( .A1(n2), .A2(n32), .B1(net106765), .B2(n10), .ZN(n80) );
  INV_X1 U64 ( .A(data_in[24]), .ZN(n32) );
  OAI22_X1 U65 ( .A1(n2), .A2(n30), .B1(net106766), .B2(n10), .ZN(n82) );
  INV_X1 U66 ( .A(data_in[25]), .ZN(n30) );
  NAND2_X1 U67 ( .A1(load), .A2(enable), .ZN(n29) );
  INV_X1 U68 ( .A(reset), .ZN(n14) );
endmodule


module Mux_NBit_2x1_NBIT_IN26 ( port0, port1, sel, portY );
  input [25:0] port0;
  input [25:0] port1;
  output [25:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, n28, n30, n31,
         n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n1;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;

  INV_X2 U1 ( .A(sel), .ZN(n1) );
  INV_X1 U2 ( .A(n44), .ZN(N2) );
  AOI22_X1 U3 ( .A1(port0[0]), .A2(n1), .B1(port1[0]), .B2(sel), .ZN(n44) );
  INV_X1 U4 ( .A(n35), .ZN(N3) );
  AOI22_X1 U5 ( .A1(port0[1]), .A2(n1), .B1(port1[1]), .B2(sel), .ZN(n35) );
  INV_X1 U6 ( .A(n34), .ZN(N4) );
  AOI22_X1 U7 ( .A1(port0[2]), .A2(n1), .B1(port1[2]), .B2(sel), .ZN(n34) );
  INV_X1 U8 ( .A(n33), .ZN(N5) );
  AOI22_X1 U9 ( .A1(port0[3]), .A2(n1), .B1(port1[3]), .B2(sel), .ZN(n33) );
  INV_X1 U10 ( .A(n32), .ZN(N6) );
  AOI22_X1 U11 ( .A1(port0[4]), .A2(n1), .B1(port1[4]), .B2(sel), .ZN(n32) );
  INV_X1 U12 ( .A(n31), .ZN(N7) );
  AOI22_X1 U13 ( .A1(port0[5]), .A2(n1), .B1(port1[5]), .B2(sel), .ZN(n31) );
  INV_X1 U14 ( .A(n30), .ZN(N8) );
  AOI22_X1 U15 ( .A1(port0[6]), .A2(n1), .B1(port1[6]), .B2(sel), .ZN(n30) );
  INV_X1 U16 ( .A(n28), .ZN(N9) );
  AOI22_X1 U17 ( .A1(port0[7]), .A2(n1), .B1(sel), .B2(port1[7]), .ZN(n28) );
  INV_X1 U18 ( .A(n54), .ZN(N10) );
  AOI22_X1 U19 ( .A1(port0[8]), .A2(n1), .B1(port1[8]), .B2(sel), .ZN(n54) );
  INV_X1 U20 ( .A(n53), .ZN(N11) );
  AOI22_X1 U21 ( .A1(port0[9]), .A2(n1), .B1(port1[9]), .B2(sel), .ZN(n53) );
  INV_X1 U22 ( .A(n52), .ZN(N12) );
  AOI22_X1 U23 ( .A1(port0[10]), .A2(n1), .B1(port1[10]), .B2(sel), .ZN(n52)
         );
  INV_X1 U24 ( .A(n51), .ZN(N13) );
  AOI22_X1 U25 ( .A1(port0[11]), .A2(n1), .B1(port1[11]), .B2(sel), .ZN(n51)
         );
  INV_X1 U26 ( .A(n50), .ZN(N14) );
  AOI22_X1 U27 ( .A1(port0[12]), .A2(n1), .B1(port1[12]), .B2(sel), .ZN(n50)
         );
  INV_X1 U28 ( .A(n49), .ZN(N15) );
  AOI22_X1 U29 ( .A1(port0[13]), .A2(n1), .B1(port1[13]), .B2(sel), .ZN(n49)
         );
  INV_X1 U30 ( .A(n48), .ZN(N16) );
  AOI22_X1 U31 ( .A1(port0[14]), .A2(n1), .B1(port1[14]), .B2(sel), .ZN(n48)
         );
  INV_X1 U32 ( .A(n47), .ZN(N17) );
  AOI22_X1 U33 ( .A1(port0[15]), .A2(n1), .B1(port1[15]), .B2(sel), .ZN(n47)
         );
  INV_X1 U34 ( .A(n46), .ZN(N18) );
  AOI22_X1 U35 ( .A1(port0[16]), .A2(n1), .B1(port1[16]), .B2(sel), .ZN(n46)
         );
  INV_X1 U36 ( .A(n45), .ZN(N19) );
  AOI22_X1 U37 ( .A1(port0[17]), .A2(n1), .B1(port1[17]), .B2(sel), .ZN(n45)
         );
  INV_X1 U38 ( .A(n43), .ZN(N20) );
  AOI22_X1 U39 ( .A1(port0[18]), .A2(n1), .B1(port1[18]), .B2(sel), .ZN(n43)
         );
  INV_X1 U40 ( .A(n42), .ZN(N21) );
  AOI22_X1 U41 ( .A1(port0[19]), .A2(n1), .B1(port1[19]), .B2(sel), .ZN(n42)
         );
  INV_X1 U42 ( .A(n41), .ZN(N22) );
  AOI22_X1 U43 ( .A1(port0[20]), .A2(n1), .B1(port1[20]), .B2(sel), .ZN(n41)
         );
  INV_X1 U44 ( .A(n40), .ZN(N23) );
  AOI22_X1 U45 ( .A1(port0[21]), .A2(n1), .B1(port1[21]), .B2(sel), .ZN(n40)
         );
  INV_X1 U46 ( .A(n39), .ZN(N24) );
  AOI22_X1 U47 ( .A1(port0[22]), .A2(n1), .B1(port1[22]), .B2(sel), .ZN(n39)
         );
  INV_X1 U48 ( .A(n38), .ZN(N25) );
  AOI22_X1 U49 ( .A1(port0[23]), .A2(n1), .B1(port1[23]), .B2(sel), .ZN(n38)
         );
  INV_X1 U50 ( .A(n37), .ZN(N26) );
  AOI22_X1 U51 ( .A1(port0[24]), .A2(n1), .B1(port1[24]), .B2(sel), .ZN(n37)
         );
  INV_X1 U52 ( .A(n36), .ZN(N27) );
  AOI22_X1 U53 ( .A1(port0[25]), .A2(n1), .B1(port1[25]), .B2(sel), .ZN(n36)
         );
endmodule


module FCU ( FCU_enable, FCU_IF_ID_Op, FCU_ID_EX_Op, FCU_EX_MEM_Op, 
        FCU_MEM_WB_Op, FCU_IF_ID_6_10, FCU_IF_ID_11_15, FCU_ID_EX_6_10, 
        FCU_ID_EX_11_15, FCU_ID_EX_16_20, FCU_EX_MEM_11_15, FCU_EX_MEM_16_20, 
        FCU_MEM_WB_11_15, FCU_MEM_WB_16_20, FCU_IF_ID_MUX, FCU_ID_EX_TOP_MUX, 
        FCU_ID_EX_BOT_MUX, FCU_EX_MEM_MUX, FCU_IF_ID_is_branch, 
        FCU_ID_EX_is_store, FCU_IF_ID_is_branch_or_jmp, FCU_IF_ID_is_jmp_r, 
        FCU_insert_stall );
  input [5:0] FCU_IF_ID_Op;
  input [5:0] FCU_ID_EX_Op;
  input [5:0] FCU_EX_MEM_Op;
  input [5:0] FCU_MEM_WB_Op;
  input [4:0] FCU_IF_ID_6_10;
  input [4:0] FCU_IF_ID_11_15;
  input [4:0] FCU_ID_EX_6_10;
  input [4:0] FCU_ID_EX_11_15;
  input [4:0] FCU_ID_EX_16_20;
  input [4:0] FCU_EX_MEM_11_15;
  input [4:0] FCU_EX_MEM_16_20;
  input [4:0] FCU_MEM_WB_11_15;
  input [4:0] FCU_MEM_WB_16_20;
  output [1:0] FCU_IF_ID_MUX;
  output [1:0] FCU_ID_EX_TOP_MUX;
  output [1:0] FCU_ID_EX_BOT_MUX;
  input FCU_enable;
  output FCU_EX_MEM_MUX, FCU_IF_ID_is_branch, FCU_ID_EX_is_store,
         FCU_IF_ID_is_branch_or_jmp, FCU_IF_ID_is_jmp_r, FCU_insert_stall;
  wire   s_stall_de, s_id_ex_is_load, s_if_id_is_reg, s_if_id_is_imm,
         s_if_id_is_load, s_if_id_is_store, s_ex_mem_is_load, s_id_ex_is_reg,
         s_id_ex_is_imm, s_ex_mem_is_reg, s_ex_mem_is_imm, s_mem_wb_is_load,
         s_stall_mem, s_stall_ex, s_mem_wb_is_reg, s_mem_wb_is_imm,
         s_ex_mem_is_store, N309, N310, N311, N312, N319, N326, N333, N340,
         N341, N343, N344, N346, N347, N349, N350, N352, N355, N358, N361,
         N364, N365, N366, N367, n241, n48, n49, n50, n51, n52, n53, n54, n55,
         n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n68, n69,
         n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83,
         n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97,
         n98, n99, n100, n101, n102, n103, n104, n105, n106, n107, n108, n109,
         n110, n111, n112, n113, n114, n115, n116, n117, n118, n119, n120,
         n121, n122, n123, n124, n125, n126, n127, n128, n129, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n148, n149, n150, n151, n152, n153,
         n154, n155, n157, n158, n159, n160, n161, n162, n163, n164, n165,
         n167, n168, n169, n170, n171, n172, n173, n174, n175, n176, n178,
         n179, n180, n181, n182, n183, n184, n185, n186, n187, n188, n189,
         n190, n191, n192, n193, n194, n195, n196, n197, n198, n199, n200,
         n201, n202, n203, n204, n205, n206, n207, n208, n210, n211, n212,
         n213, n214, n215, n217, n220, n221, n222, n223, n224, n225, n226,
         n227, n228, n229, n230, n231, n232, n233, n234, n235, n236, n237,
         n238, n243, n244, n245, n249, n250, n251, n252, n254, n255, n258,
         n259, n263, n264, n265, n266, n267, n268, n269, n270, n271, n272,
         n273, n274, n275, n276, n277, n278, n279, n280, n281, n242, n246,
         n247, n248, n253, n256, n257, n260, n261, n262, n282, n283, n284,
         n285, n286, n287, n289, n290, n291, n292, n293, n294, n295, n296,
         n297, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n317, n318,
         n319, n320, n321, n322, n323, n324, n325, n326, n327, n328;
  assign FCU_insert_stall = s_stall_de;
  assign N341 = FCU_IF_ID_Op[5];
  assign N344 = FCU_ID_EX_Op[5];
  assign N347 = FCU_EX_MEM_Op[5];
  assign N350 = FCU_MEM_WB_Op[5];

  DLH_X1 FCU_IF_ID_is_branch_reg ( .G(n326), .D(N366), .Q(FCU_IF_ID_is_branch)
         );
  DLH_X1 s_if_id_is_reg_reg ( .G(n326), .D(N309), .Q(s_if_id_is_reg) );
  DLH_X1 s_id_ex_is_reg_reg ( .G(n326), .D(N310), .Q(s_id_ex_is_reg) );
  DLH_X1 s_ex_mem_is_reg_reg ( .G(n326), .D(N311), .Q(s_ex_mem_is_reg) );
  DLH_X1 s_mem_wb_is_reg_reg ( .G(n326), .D(N312), .Q(s_mem_wb_is_reg) );
  DLH_X1 s_if_id_is_imm_reg ( .G(n326), .D(N319), .Q(s_if_id_is_imm) );
  DLH_X1 s_id_ex_is_imm_reg ( .G(n326), .D(N326), .Q(s_id_ex_is_imm) );
  DLH_X1 s_ex_mem_is_imm_reg ( .G(n326), .D(N333), .Q(s_ex_mem_is_imm) );
  DLH_X1 s_mem_wb_is_imm_reg ( .G(n326), .D(N340), .Q(s_mem_wb_is_imm) );
  DLH_X1 s_if_id_is_load_reg ( .G(n326), .D(N343), .Q(s_if_id_is_load) );
  DLH_X1 s_id_ex_is_load_reg ( .G(n326), .D(N346), .Q(s_id_ex_is_load) );
  DLH_X1 s_ex_mem_is_load_reg ( .G(n326), .D(N349), .Q(s_ex_mem_is_load) );
  DLH_X1 s_mem_wb_is_load_reg ( .G(n326), .D(N352), .Q(s_mem_wb_is_load) );
  DLH_X1 s_if_id_is_store_reg ( .G(n326), .D(N355), .Q(s_if_id_is_store) );
  DLH_X1 s_id_ex_is_store_reg ( .G(n326), .D(N358), .Q(FCU_ID_EX_is_store) );
  DLH_X1 s_ex_mem_is_store_reg ( .G(n326), .D(N361), .Q(s_ex_mem_is_store) );
  DLH_X1 s_if_id_is_jmp_r_reg ( .G(N367), .D(N364), .Q(FCU_IF_ID_is_jmp_r) );
  DLH_X1 s_if_id_is_jmp_reg ( .G(n326), .D(N365), .Q(
        FCU_IF_ID_is_branch_or_jmp) );
  DLH_X1 s_stall_ex_reg ( .G(n326), .D(n241), .Q(s_stall_ex) );
  DLH_X1 s_stall_mem_reg ( .G(n326), .D(s_stall_ex), .Q(s_stall_mem) );
  NAND3_X1 U233 ( .A1(n52), .A2(n53), .A3(s_id_ex_is_load), .ZN(n51) );
  XOR2_X1 U234 ( .A(FCU_IF_ID_11_15[4]), .B(FCU_ID_EX_11_15[4]), .Z(n63) );
  XOR2_X1 U235 ( .A(FCU_IF_ID_11_15[3]), .B(FCU_ID_EX_11_15[3]), .Z(n62) );
  NAND3_X1 U236 ( .A1(n64), .A2(n65), .A3(n66), .ZN(n61) );
  XOR2_X1 U237 ( .A(FCU_IF_ID_6_10[3]), .B(FCU_ID_EX_11_15[3]), .Z(n78) );
  XOR2_X1 U238 ( .A(FCU_IF_ID_6_10[1]), .B(FCU_ID_EX_16_20[1]), .Z(n84) );
  XOR2_X1 U239 ( .A(FCU_IF_ID_6_10[3]), .B(FCU_ID_EX_16_20[3]), .Z(n88) );
  XOR2_X1 U240 ( .A(FCU_IF_ID_6_10[0]), .B(FCU_ID_EX_16_20[0]), .Z(n87) );
  XOR2_X1 U241 ( .A(FCU_IF_ID_6_10[2]), .B(FCU_ID_EX_16_20[2]), .Z(n86) );
  NAND3_X1 U242 ( .A1(N347), .A2(n121), .A3(FCU_EX_MEM_Op[4]), .ZN(n120) );
  NAND3_X1 U243 ( .A1(N344), .A2(n129), .A3(FCU_ID_EX_Op[4]), .ZN(n128) );
  NAND3_X1 U244 ( .A1(N341), .A2(n137), .A3(FCU_IF_ID_Op[4]), .ZN(n136) );
  NAND3_X1 U245 ( .A1(FCU_IF_ID_is_branch_or_jmp), .A2(n53), .A3(n326), .ZN(
        n146) );
  XOR2_X1 U246 ( .A(FCU_IF_ID_6_10[3]), .B(FCU_EX_MEM_16_20[3]), .Z(n161) );
  NAND3_X1 U247 ( .A1(n165), .A2(n321), .A3(n167), .ZN(n160) );
  XOR2_X1 U248 ( .A(FCU_MEM_WB_11_15[1]), .B(FCU_IF_ID_6_10[1]), .Z(n150) );
  XOR2_X1 U249 ( .A(FCU_MEM_WB_11_15[0]), .B(FCU_IF_ID_6_10[0]), .Z(n152) );
  XOR2_X1 U250 ( .A(FCU_MEM_WB_11_15[3]), .B(FCU_IF_ID_6_10[3]), .Z(n147) );
  XOR2_X1 U251 ( .A(FCU_ID_EX_6_10[2]), .B(FCU_EX_MEM_16_20[2]), .Z(n212) );
  XOR2_X1 U252 ( .A(FCU_ID_EX_6_10[3]), .B(FCU_EX_MEM_16_20[3]), .Z(n211) );
  XOR2_X1 U253 ( .A(FCU_ID_EX_6_10[4]), .B(FCU_EX_MEM_16_20[4]), .Z(n210) );
  NAND3_X1 U256 ( .A1(n220), .A2(n221), .A3(n222), .ZN(n215) );
  NAND3_X1 U259 ( .A1(n157), .A2(n249), .A3(n250), .ZN(n245) );
  XOR2_X1 U261 ( .A(FCU_ID_EX_11_15[3]), .B(FCU_EX_MEM_16_20[3]), .Z(n255) );
  NAND3_X1 U263 ( .A1(n194), .A2(n193), .A3(n192), .ZN(n272) );
  NOR2_X1 U3 ( .A1(n327), .A2(n178), .ZN(n242) );
  INV_X1 U4 ( .A(n328), .ZN(n326) );
  CLKBUF_X1 U5 ( .A(FCU_EX_MEM_16_20[1]), .Z(n246) );
  AOI21_X1 U6 ( .B1(n296), .B2(n297), .A(n295), .ZN(n247) );
  BUF_X1 U7 ( .A(FCU_EX_MEM_11_15[4]), .Z(n248) );
  AND3_X2 U8 ( .A1(n291), .A2(n292), .A3(n293), .ZN(n243) );
  INV_X1 U9 ( .A(s_ex_mem_is_reg), .ZN(n295) );
  OR3_X1 U10 ( .A1(FCU_EX_MEM_11_15[3]), .A2(FCU_EX_MEM_11_15[4]), .A3(
        FCU_EX_MEM_11_15[2]), .ZN(n251) );
  BUF_X1 U11 ( .A(FCU_ID_EX_6_10[2]), .Z(n305) );
  OR2_X1 U12 ( .A1(n224), .A2(n225), .ZN(n253) );
  OR2_X1 U13 ( .A1(n223), .A2(n225), .ZN(n256) );
  OAI21_X1 U14 ( .B1(n318), .B2(n309), .A(s_ex_mem_is_imm), .ZN(n257) );
  XNOR2_X1 U15 ( .A(FCU_ID_EX_6_10[1]), .B(FCU_EX_MEM_11_15[1]), .ZN(n260) );
  AND3_X1 U16 ( .A1(n261), .A2(n262), .A3(n282), .ZN(n238) );
  XOR2_X1 U17 ( .A(n198), .B(FCU_ID_EX_11_15[0]), .Z(n261) );
  XOR2_X1 U18 ( .A(n199), .B(FCU_ID_EX_11_15[1]), .Z(n262) );
  XOR2_X1 U19 ( .A(n176), .B(FCU_ID_EX_11_15[2]), .Z(n282) );
  CLKBUF_X1 U20 ( .A(FCU_ID_EX_6_10[4]), .Z(n283) );
  BUF_X1 U21 ( .A(FCU_EX_MEM_11_15[2]), .Z(n284) );
  CLKBUF_X1 U22 ( .A(FCU_ID_EX_11_15[1]), .Z(n285) );
  XNOR2_X1 U23 ( .A(FCU_ID_EX_6_10[0]), .B(FCU_EX_MEM_11_15[0]), .ZN(n286) );
  NOR3_X1 U24 ( .A1(n257), .A2(n215), .A3(n310), .ZN(n287) );
  NAND2_X1 U25 ( .A1(n289), .A2(n290), .ZN(FCU_ID_EX_BOT_MUX[1]) );
  OR2_X1 U26 ( .A1(n226), .A2(n253), .ZN(n289) );
  OR2_X1 U27 ( .A1(n226), .A2(n256), .ZN(n290) );
  AND3_X1 U28 ( .A1(n294), .A2(n258), .A3(n259), .ZN(n291) );
  XNOR2_X1 U29 ( .A(n308), .B(FCU_ID_EX_11_15[2]), .ZN(n292) );
  NOR2_X1 U30 ( .A1(n255), .A2(n254), .ZN(n293) );
  AOI21_X1 U31 ( .B1(n296), .B2(n297), .A(n295), .ZN(n294) );
  NOR3_X1 U32 ( .A1(FCU_EX_MEM_16_20[3]), .A2(FCU_EX_MEM_16_20[2]), .A3(
        FCU_EX_MEM_16_20[4]), .ZN(n296) );
  NOR2_X1 U33 ( .A1(FCU_EX_MEM_16_20[1]), .A2(FCU_EX_MEM_16_20[0]), .ZN(n297)
         );
  AND4_X1 U34 ( .A1(n324), .A2(n214), .A3(n213), .A4(n247), .ZN(n208) );
  NAND2_X1 U35 ( .A1(n260), .A2(n286), .ZN(n310) );
  AND2_X1 U36 ( .A1(n205), .A2(n313), .ZN(FCU_ID_EX_TOP_MUX[1]) );
  OAI211_X1 U37 ( .C1(n207), .C2(n208), .A(s_stall_mem), .B(n242), .ZN(n298)
         );
  INV_X1 U38 ( .A(n298), .ZN(FCU_ID_EX_TOP_MUX[0]) );
  OAI211_X1 U39 ( .C1(n243), .C2(n244), .A(s_stall_mem), .B(n323), .ZN(n299)
         );
  INV_X1 U40 ( .A(n299), .ZN(FCU_ID_EX_BOT_MUX[0]) );
  CLKBUF_X1 U41 ( .A(FCU_EX_MEM_11_15[0]), .Z(n300) );
  NAND3_X1 U42 ( .A1(n302), .A2(n303), .A3(n304), .ZN(n301) );
  XNOR2_X1 U43 ( .A(n248), .B(FCU_ID_EX_11_15[4]), .ZN(n302) );
  XNOR2_X1 U44 ( .A(FCU_ID_EX_11_15[1]), .B(FCU_EX_MEM_11_15[1]), .ZN(n303) );
  XNOR2_X1 U45 ( .A(n284), .B(FCU_ID_EX_11_15[2]), .ZN(n304) );
  CLKBUF_X1 U46 ( .A(FCU_EX_MEM_16_20[4]), .Z(n306) );
  BUF_X1 U47 ( .A(FCU_EX_MEM_16_20[0]), .Z(n307) );
  CLKBUF_X1 U48 ( .A(FCU_EX_MEM_16_20[2]), .Z(n308) );
  OR3_X1 U49 ( .A1(FCU_EX_MEM_11_15[3]), .A2(FCU_EX_MEM_11_15[2]), .A3(
        FCU_EX_MEM_11_15[4]), .ZN(n309) );
  CLKBUF_X1 U50 ( .A(n284), .Z(n311) );
  CLKBUF_X1 U51 ( .A(FCU_ID_EX_11_15[2]), .Z(n312) );
  NOR3_X1 U52 ( .A1(n179), .A2(n328), .A3(n178), .ZN(n313) );
  CLKBUF_X1 U53 ( .A(n308), .Z(n314) );
  CLKBUF_X1 U54 ( .A(n157), .Z(n315) );
  CLKBUF_X1 U55 ( .A(FCU_EX_MEM_11_15[1]), .Z(n316) );
  CLKBUF_X1 U56 ( .A(FCU_ID_EX_11_15[0]), .Z(n317) );
  BUF_X1 U57 ( .A(n252), .Z(n318) );
  CLKBUF_X1 U58 ( .A(FCU_EX_MEM_11_15[3]), .Z(n319) );
  CLKBUF_X1 U59 ( .A(n248), .Z(n320) );
  CLKBUF_X1 U60 ( .A(n294), .Z(n321) );
  XOR2_X1 U61 ( .A(FCU_ID_EX_11_15[0]), .B(FCU_EX_MEM_16_20[0]), .Z(n254) );
  NOR3_X1 U62 ( .A1(n322), .A2(n215), .A3(n310), .ZN(n207) );
  OAI21_X1 U63 ( .B1(n318), .B2(n309), .A(s_ex_mem_is_imm), .ZN(n322) );
  NOR2_X1 U64 ( .A1(n328), .A2(n83), .ZN(n323) );
  NOR3_X1 U65 ( .A1(n211), .A2(n210), .A3(n212), .ZN(n324) );
  NOR2_X1 U66 ( .A1(n245), .A2(n301), .ZN(n244) );
  INV_X1 U67 ( .A(FCU_enable), .ZN(n328) );
  AND2_X1 U68 ( .A1(N365), .A2(n326), .ZN(N367) );
  AOI22_X1 U69 ( .A1(n181), .A2(n180), .B1(n182), .B2(n183), .ZN(n179) );
  NOR3_X1 U70 ( .A1(n189), .A2(n190), .A3(n191), .ZN(n182) );
  INV_X1 U71 ( .A(n196), .ZN(n236) );
  INV_X1 U72 ( .A(n185), .ZN(n229) );
  NOR2_X1 U73 ( .A1(n89), .A2(n90), .ZN(n67) );
  INV_X1 U74 ( .A(n89), .ZN(n53) );
  NAND2_X1 U75 ( .A1(n326), .A2(n48), .ZN(s_stall_de) );
  INV_X1 U76 ( .A(n55), .ZN(n57) );
  NOR4_X1 U77 ( .A1(n154), .A2(n155), .A3(n50), .A4(n328), .ZN(
        FCU_IF_ID_MUX[0]) );
  NOR4_X1 U78 ( .A1(n175), .A2(n151), .A3(n152), .A4(n150), .ZN(n154) );
  OR3_X1 U79 ( .A1(n148), .A2(n147), .A3(n153), .ZN(n175) );
  INV_X1 U80 ( .A(n90), .ZN(n158) );
  NOR2_X1 U81 ( .A1(n113), .A2(n114), .ZN(n102) );
  AOI21_X1 U82 ( .B1(n113), .B2(n114), .A(n115), .ZN(n111) );
  OAI21_X1 U83 ( .B1(n92), .B2(n93), .A(n91), .ZN(N365) );
  NOR2_X1 U84 ( .A1(n97), .A2(n98), .ZN(N361) );
  NOR2_X1 U85 ( .A1(n99), .A2(n100), .ZN(N358) );
  INV_X1 U86 ( .A(n91), .ZN(N366) );
  INV_X1 U87 ( .A(n48), .ZN(n241) );
  NAND2_X1 U88 ( .A1(FCU_enable), .A2(s_id_ex_is_reg), .ZN(n225) );
  NAND4_X1 U89 ( .A1(n235), .A2(n236), .A3(n237), .A4(n238), .ZN(n223) );
  NAND4_X1 U90 ( .A1(n228), .A2(n229), .A3(n230), .A4(n231), .ZN(n224) );
  NOR3_X1 U91 ( .A1(n232), .A2(n233), .A3(n234), .ZN(n231) );
  XNOR2_X1 U92 ( .A(n192), .B(FCU_ID_EX_11_15[2]), .ZN(n234) );
  NOR3_X1 U93 ( .A1(n196), .A2(n195), .A3(n197), .ZN(n181) );
  XNOR2_X1 U94 ( .A(n199), .B(FCU_ID_EX_6_10[1]), .ZN(n195) );
  XNOR2_X1 U95 ( .A(n198), .B(FCU_ID_EX_6_10[0]), .ZN(n197) );
  NOR3_X1 U96 ( .A1(n184), .A2(n185), .A3(n186), .ZN(n183) );
  XNOR2_X1 U97 ( .A(n188), .B(FCU_ID_EX_6_10[0]), .ZN(n184) );
  XNOR2_X1 U98 ( .A(n187), .B(FCU_ID_EX_6_10[1]), .ZN(n186) );
  NOR3_X1 U99 ( .A1(n200), .A2(n201), .A3(n202), .ZN(n180) );
  XNOR2_X1 U100 ( .A(n176), .B(n305), .ZN(n201) );
  XNOR2_X1 U101 ( .A(n204), .B(n283), .ZN(n200) );
  XNOR2_X1 U102 ( .A(n203), .B(FCU_ID_EX_6_10[3]), .ZN(n202) );
  OAI21_X1 U103 ( .B1(n272), .B2(n273), .A(s_mem_wb_is_reg), .ZN(n185) );
  NAND2_X1 U104 ( .A1(n188), .A2(n187), .ZN(n273) );
  OAI21_X1 U105 ( .B1(s_mem_wb_is_load), .B2(s_mem_wb_is_imm), .A(n280), .ZN(
        n196) );
  NAND4_X1 U106 ( .A1(n203), .A2(n204), .A3(n176), .A4(n281), .ZN(n280) );
  NOR2_X1 U107 ( .A1(FCU_MEM_WB_11_15[1]), .A2(FCU_MEM_WB_11_15[0]), .ZN(n281)
         );
  INV_X1 U108 ( .A(FCU_MEM_WB_11_15[2]), .ZN(n176) );
  XNOR2_X1 U109 ( .A(FCU_MEM_WB_16_20[3]), .B(FCU_ID_EX_11_15[3]), .ZN(n230)
         );
  XNOR2_X1 U110 ( .A(FCU_MEM_WB_11_15[3]), .B(FCU_ID_EX_11_15[3]), .ZN(n237)
         );
  XNOR2_X1 U111 ( .A(n192), .B(n305), .ZN(n191) );
  XNOR2_X1 U112 ( .A(n193), .B(FCU_ID_EX_6_10[4]), .ZN(n190) );
  XNOR2_X1 U113 ( .A(FCU_ID_EX_6_10[3]), .B(n194), .ZN(n189) );
  INV_X1 U114 ( .A(FCU_MEM_WB_16_20[2]), .ZN(n192) );
  INV_X1 U115 ( .A(FCU_MEM_WB_16_20[1]), .ZN(n187) );
  INV_X1 U116 ( .A(FCU_MEM_WB_11_15[4]), .ZN(n204) );
  INV_X1 U117 ( .A(FCU_MEM_WB_11_15[3]), .ZN(n203) );
  INV_X1 U118 ( .A(FCU_MEM_WB_16_20[0]), .ZN(n188) );
  INV_X1 U119 ( .A(FCU_MEM_WB_16_20[3]), .ZN(n194) );
  INV_X1 U120 ( .A(FCU_MEM_WB_16_20[4]), .ZN(n193) );
  INV_X1 U121 ( .A(FCU_MEM_WB_11_15[0]), .ZN(n198) );
  INV_X1 U122 ( .A(FCU_MEM_WB_11_15[1]), .ZN(n199) );
  NOR4_X1 U123 ( .A1(FCU_IF_ID_6_10[3]), .A2(FCU_IF_ID_6_10[4]), .A3(
        FCU_IF_ID_6_10[2]), .A4(n149), .ZN(n89) );
  OR2_X1 U124 ( .A1(FCU_IF_ID_6_10[1]), .A2(FCU_IF_ID_6_10[0]), .ZN(n149) );
  NAND4_X1 U125 ( .A1(n74), .A2(n75), .A3(n76), .A4(n77), .ZN(n55) );
  XNOR2_X1 U126 ( .A(n312), .B(FCU_IF_ID_6_10[2]), .ZN(n76) );
  NOR3_X1 U127 ( .A1(n55), .A2(n71), .A3(n72), .ZN(n70) );
  NOR3_X1 U128 ( .A1(n61), .A2(n62), .A3(n63), .ZN(n58) );
  OAI21_X1 U129 ( .B1(n49), .B2(n50), .A(n51), .ZN(n48) );
  AOI221_X1 U130 ( .B1(n67), .B2(s_ex_mem_is_load), .C1(n68), .C2(n69), .A(n70), .ZN(n49) );
  NOR3_X1 U131 ( .A1(n86), .A2(n87), .A3(n88), .ZN(n68) );
  INV_X1 U132 ( .A(FCU_IF_ID_6_10[4]), .ZN(n80) );
  NAND4_X1 U133 ( .A1(n168), .A2(n169), .A3(n170), .A4(n171), .ZN(n90) );
  XNOR2_X1 U134 ( .A(n325), .B(FCU_IF_ID_6_10[0]), .ZN(n169) );
  NOR4_X1 U135 ( .A1(n81), .A2(n82), .A3(n83), .A4(n84), .ZN(n69) );
  AND2_X1 U136 ( .A1(n80), .A2(FCU_ID_EX_16_20[4]), .ZN(n82) );
  AOI21_X1 U137 ( .B1(n80), .B2(n85), .A(FCU_ID_EX_16_20[4]), .ZN(n81) );
  XNOR2_X1 U138 ( .A(FCU_IF_ID_11_15[2]), .B(n312), .ZN(n65) );
  NOR2_X1 U139 ( .A1(n78), .A2(n79), .ZN(n77) );
  NOR2_X1 U140 ( .A1(n172), .A2(n173), .ZN(n171) );
  XNOR2_X1 U141 ( .A(FCU_IF_ID_6_10[2]), .B(n174), .ZN(n172) );
  OR4_X1 U142 ( .A1(FCU_ID_EX_16_20[0]), .A2(FCU_ID_EX_16_20[1]), .A3(
        FCU_ID_EX_16_20[2]), .A4(FCU_ID_EX_16_20[3]), .ZN(n85) );
  OAI21_X1 U143 ( .B1(n54), .B2(n55), .A(n56), .ZN(n52) );
  NOR4_X1 U144 ( .A1(s_if_id_is_store), .A2(s_if_id_is_load), .A3(
        s_if_id_is_imm), .A4(FCU_IF_ID_is_branch_or_jmp), .ZN(n54) );
  OAI211_X1 U145 ( .C1(n57), .C2(n58), .A(n59), .B(s_if_id_is_reg), .ZN(n56)
         );
  OR4_X1 U146 ( .A1(FCU_IF_ID_11_15[3]), .A2(FCU_IF_ID_11_15[4]), .A3(
        FCU_IF_ID_11_15[2]), .A4(n60), .ZN(n59) );
  OR2_X1 U147 ( .A1(FCU_IF_ID_11_15[1]), .A2(FCU_IF_ID_11_15[0]), .ZN(n60) );
  NOR4_X1 U148 ( .A1(n145), .A2(n146), .A3(n147), .A4(n148), .ZN(
        FCU_IF_ID_MUX[1]) );
  OR4_X1 U149 ( .A1(n150), .A2(n151), .A3(n152), .A4(n153), .ZN(n145) );
  NOR4_X1 U150 ( .A1(n160), .A2(n161), .A3(n162), .A4(n163), .ZN(n159) );
  XNOR2_X1 U151 ( .A(FCU_MEM_WB_11_15[4]), .B(n80), .ZN(n148) );
  XNOR2_X1 U152 ( .A(n176), .B(FCU_IF_ID_6_10[2]), .ZN(n153) );
  AOI211_X1 U153 ( .C1(n263), .C2(n264), .A(n265), .B(n328), .ZN(
        FCU_EX_MEM_MUX) );
  INV_X1 U154 ( .A(s_ex_mem_is_store), .ZN(n265) );
  NAND4_X1 U155 ( .A1(n274), .A2(n236), .A3(n275), .A4(n276), .ZN(n263) );
  NAND4_X1 U156 ( .A1(n266), .A2(n229), .A3(n267), .A4(n268), .ZN(n264) );
  INV_X1 U157 ( .A(n72), .ZN(n206) );
  NOR3_X1 U158 ( .A1(FCU_MEM_WB_Op[2]), .A2(FCU_MEM_WB_Op[3]), .A3(
        FCU_MEM_WB_Op[1]), .ZN(n112) );
  AOI211_X1 U159 ( .C1(FCU_EX_MEM_Op[0]), .C2(n125), .A(n126), .B(
        FCU_EX_MEM_Op[3]), .ZN(n123) );
  INV_X1 U160 ( .A(FCU_EX_MEM_Op[1]), .ZN(n125) );
  NAND2_X1 U161 ( .A1(FCU_EX_MEM_Op[4]), .A2(FCU_EX_MEM_Op[2]), .ZN(n126) );
  AOI211_X1 U162 ( .C1(FCU_ID_EX_Op[0]), .C2(n133), .A(n134), .B(
        FCU_ID_EX_Op[3]), .ZN(n131) );
  INV_X1 U163 ( .A(FCU_ID_EX_Op[1]), .ZN(n133) );
  NAND2_X1 U164 ( .A1(FCU_ID_EX_Op[4]), .A2(FCU_ID_EX_Op[2]), .ZN(n134) );
  AOI211_X1 U165 ( .C1(FCU_IF_ID_Op[0]), .C2(n93), .A(n141), .B(
        FCU_IF_ID_Op[3]), .ZN(n139) );
  NAND2_X1 U166 ( .A1(FCU_IF_ID_Op[4]), .A2(FCU_IF_ID_Op[2]), .ZN(n141) );
  AOI211_X1 U167 ( .C1(FCU_MEM_WB_Op[0]), .C2(n114), .A(n118), .B(
        FCU_MEM_WB_Op[3]), .ZN(n116) );
  NAND2_X1 U168 ( .A1(FCU_MEM_WB_Op[4]), .A2(FCU_MEM_WB_Op[2]), .ZN(n118) );
  NOR4_X1 U169 ( .A1(FCU_IF_ID_Op[4]), .A2(FCU_IF_ID_Op[2]), .A3(n95), .A4(
        n101), .ZN(N355) );
  NOR4_X1 U170 ( .A1(FCU_EX_MEM_Op[4]), .A2(FCU_EX_MEM_Op[3]), .A3(n104), .A4(
        n105), .ZN(N349) );
  NOR4_X1 U171 ( .A1(FCU_ID_EX_Op[4]), .A2(FCU_ID_EX_Op[3]), .A3(n106), .A4(
        n107), .ZN(N346) );
  NOR4_X1 U172 ( .A1(FCU_IF_ID_Op[4]), .A2(FCU_IF_ID_Op[3]), .A3(n108), .A4(
        n101), .ZN(N343) );
  NOR4_X1 U173 ( .A1(FCU_MEM_WB_Op[4]), .A2(FCU_MEM_WB_Op[3]), .A3(n102), .A4(
        n103), .ZN(N352) );
  NOR3_X1 U174 ( .A1(n269), .A2(n270), .A3(n271), .ZN(n268) );
  NOR3_X1 U175 ( .A1(n277), .A2(n278), .A3(n279), .ZN(n276) );
  NAND4_X1 U176 ( .A1(FCU_IF_ID_Op[2]), .A2(n93), .A3(n94), .A4(n95), .ZN(n91)
         );
  NOR2_X1 U177 ( .A1(N341), .A2(FCU_IF_ID_Op[4]), .ZN(n94) );
  NOR2_X1 U178 ( .A1(FCU_ID_EX_is_store), .A2(s_id_ex_is_imm), .ZN(n72) );
  AOI21_X1 U179 ( .B1(n104), .B2(FCU_EX_MEM_Op[4]), .A(n97), .ZN(n124) );
  AOI21_X1 U180 ( .B1(n106), .B2(FCU_ID_EX_Op[4]), .A(n99), .ZN(n132) );
  INV_X1 U181 ( .A(FCU_IF_ID_Op[3]), .ZN(n95) );
  NOR3_X1 U182 ( .A1(n92), .A2(FCU_IF_ID_Op[4]), .A3(FCU_IF_ID_Op[1]), .ZN(
        N309) );
  NOR3_X1 U183 ( .A1(n98), .A2(FCU_EX_MEM_Op[3]), .A3(FCU_EX_MEM_Op[1]), .ZN(
        N311) );
  NOR3_X1 U184 ( .A1(n100), .A2(FCU_ID_EX_Op[3]), .A3(FCU_ID_EX_Op[1]), .ZN(
        N310) );
  INV_X1 U185 ( .A(FCU_IF_ID_Op[1]), .ZN(n93) );
  NOR2_X1 U186 ( .A1(FCU_EX_MEM_Op[1]), .A2(FCU_EX_MEM_Op[2]), .ZN(n122) );
  NOR2_X1 U187 ( .A1(FCU_ID_EX_Op[1]), .A2(FCU_ID_EX_Op[2]), .ZN(n130) );
  NOR3_X1 U188 ( .A1(n142), .A2(N350), .A3(FCU_MEM_WB_Op[4]), .ZN(N312) );
  INV_X1 U189 ( .A(n112), .ZN(n142) );
  NOR3_X1 U190 ( .A1(n96), .A2(n92), .A3(n93), .ZN(N364) );
  INV_X1 U191 ( .A(FCU_IF_ID_Op[0]), .ZN(n96) );
  INV_X1 U192 ( .A(FCU_EX_MEM_Op[3]), .ZN(n97) );
  INV_X1 U193 ( .A(FCU_ID_EX_Op[3]), .ZN(n99) );
  INV_X1 U194 ( .A(N341), .ZN(n101) );
  INV_X1 U195 ( .A(N347), .ZN(n105) );
  INV_X1 U196 ( .A(N344), .ZN(n107) );
  INV_X1 U197 ( .A(FCU_MEM_WB_Op[1]), .ZN(n114) );
  XNOR2_X1 U198 ( .A(n95), .B(n138), .ZN(n137) );
  NOR2_X1 U199 ( .A1(FCU_IF_ID_Op[1]), .A2(FCU_IF_ID_Op[2]), .ZN(n138) );
  INV_X1 U200 ( .A(FCU_IF_ID_is_branch_or_jmp), .ZN(n50) );
  AND2_X1 U201 ( .A1(FCU_IF_ID_Op[2]), .A2(FCU_IF_ID_Op[1]), .ZN(n108) );
  OR3_X1 U202 ( .A1(FCU_IF_ID_Op[3]), .A2(N341), .A3(FCU_IF_ID_Op[2]), .ZN(n92) );
  AND2_X1 U203 ( .A1(FCU_EX_MEM_Op[2]), .A2(FCU_EX_MEM_Op[1]), .ZN(n104) );
  AND2_X1 U204 ( .A1(FCU_ID_EX_Op[2]), .A2(FCU_ID_EX_Op[1]), .ZN(n106) );
  OR3_X1 U205 ( .A1(FCU_EX_MEM_Op[2]), .A2(FCU_EX_MEM_Op[4]), .A3(n143), .ZN(
        n98) );
  XNOR2_X1 U206 ( .A(n105), .B(FCU_EX_MEM_Op[3]), .ZN(n143) );
  OR3_X1 U207 ( .A1(FCU_ID_EX_Op[2]), .A2(FCU_ID_EX_Op[4]), .A3(n144), .ZN(
        n100) );
  XNOR2_X1 U208 ( .A(n107), .B(FCU_ID_EX_Op[3]), .ZN(n144) );
  INV_X1 U209 ( .A(FCU_MEM_WB_Op[3]), .ZN(n115) );
  INV_X1 U210 ( .A(N350), .ZN(n103) );
  INV_X1 U211 ( .A(FCU_MEM_WB_Op[2]), .ZN(n113) );
  INV_X1 U212 ( .A(s_id_ex_is_reg), .ZN(n83) );
  INV_X1 U213 ( .A(s_mem_wb_is_load), .ZN(n151) );
  NAND2_X1 U214 ( .A1(n135), .A2(n136), .ZN(N319) );
  OAI21_X1 U215 ( .B1(n139), .B2(n140), .A(n101), .ZN(n135) );
  AOI21_X1 U216 ( .B1(n108), .B2(FCU_IF_ID_Op[4]), .A(n95), .ZN(n140) );
  NAND2_X1 U217 ( .A1(n109), .A2(n110), .ZN(N340) );
  OAI21_X1 U218 ( .B1(n116), .B2(n117), .A(n103), .ZN(n109) );
  OAI211_X1 U219 ( .C1(n111), .C2(n112), .A(N350), .B(FCU_MEM_WB_Op[4]), .ZN(
        n110) );
  AOI21_X1 U220 ( .B1(n102), .B2(FCU_MEM_WB_Op[4]), .A(n115), .ZN(n117) );
  NAND2_X1 U221 ( .A1(n119), .A2(n120), .ZN(N333) );
  OAI21_X1 U222 ( .B1(n123), .B2(n124), .A(n105), .ZN(n119) );
  XNOR2_X1 U223 ( .A(n97), .B(n122), .ZN(n121) );
  NAND2_X1 U224 ( .A1(n127), .A2(n128), .ZN(N326) );
  OAI21_X1 U225 ( .B1(n131), .B2(n132), .A(n107), .ZN(n127) );
  XNOR2_X1 U226 ( .A(n99), .B(n130), .ZN(n129) );
  XNOR2_X1 U227 ( .A(FCU_IF_ID_11_15[1]), .B(n285), .ZN(n66) );
  XNOR2_X1 U228 ( .A(n285), .B(FCU_IF_ID_6_10[1]), .ZN(n75) );
  XNOR2_X1 U229 ( .A(n187), .B(FCU_ID_EX_11_15[1]), .ZN(n233) );
  XNOR2_X1 U230 ( .A(n314), .B(FCU_IF_ID_6_10[2]), .ZN(n167) );
  XNOR2_X1 U231 ( .A(n80), .B(n306), .ZN(n163) );
  CLKBUF_X1 U232 ( .A(n300), .Z(n325) );
  NOR3_X1 U254 ( .A1(s_id_ex_is_load), .A2(s_id_ex_is_reg), .A3(n206), .ZN(
        n178) );
  INV_X1 U255 ( .A(FCU_enable), .ZN(n327) );
  AOI21_X1 U257 ( .B1(n315), .B2(n158), .A(n159), .ZN(n155) );
  XNOR2_X1 U258 ( .A(FCU_IF_ID_6_10[1]), .B(n164), .ZN(n162) );
  INV_X1 U260 ( .A(n217), .ZN(n157) );
  OR3_X1 U262 ( .A1(FCU_ID_EX_11_15[3]), .A2(FCU_ID_EX_11_15[4]), .A3(n312), 
        .ZN(n73) );
  XNOR2_X1 U264 ( .A(n80), .B(FCU_ID_EX_11_15[4]), .ZN(n79) );
  XNOR2_X1 U265 ( .A(FCU_MEM_WB_11_15[4]), .B(FCU_ID_EX_11_15[4]), .ZN(n235)
         );
  XNOR2_X1 U266 ( .A(FCU_MEM_WB_16_20[4]), .B(FCU_ID_EX_11_15[4]), .ZN(n228)
         );
  XNOR2_X1 U267 ( .A(FCU_EX_MEM_16_20[4]), .B(FCU_ID_EX_11_15[4]), .ZN(n258)
         );
  OAI21_X1 U268 ( .B1(n251), .B2(n252), .A(s_ex_mem_is_imm), .ZN(n217) );
  NOR3_X1 U269 ( .A1(n73), .A2(n285), .A3(n317), .ZN(n71) );
  XNOR2_X1 U270 ( .A(FCU_IF_ID_11_15[0]), .B(n317), .ZN(n64) );
  XNOR2_X1 U271 ( .A(n317), .B(FCU_IF_ID_6_10[0]), .ZN(n74) );
  XNOR2_X1 U272 ( .A(n188), .B(FCU_ID_EX_11_15[0]), .ZN(n232) );
  XNOR2_X1 U273 ( .A(n300), .B(FCU_ID_EX_11_15[0]), .ZN(n249) );
  XNOR2_X1 U274 ( .A(FCU_MEM_WB_16_20[0]), .B(n325), .ZN(n266) );
  XNOR2_X1 U275 ( .A(FCU_MEM_WB_11_15[0]), .B(n325), .ZN(n274) );
  XNOR2_X1 U276 ( .A(n192), .B(n311), .ZN(n270) );
  XNOR2_X1 U277 ( .A(n176), .B(n311), .ZN(n278) );
  XNOR2_X1 U278 ( .A(FCU_EX_MEM_11_15[2]), .B(FCU_ID_EX_6_10[2]), .ZN(n220) );
  INV_X1 U279 ( .A(n311), .ZN(n174) );
  XNOR2_X1 U280 ( .A(FCU_MEM_WB_16_20[1]), .B(n316), .ZN(n267) );
  XNOR2_X1 U281 ( .A(FCU_MEM_WB_11_15[1]), .B(n316), .ZN(n275) );
  XNOR2_X1 U282 ( .A(n316), .B(FCU_IF_ID_6_10[1]), .ZN(n168) );
  OR2_X1 U283 ( .A1(FCU_EX_MEM_11_15[1]), .A2(FCU_EX_MEM_11_15[0]), .ZN(n252)
         );
  XNOR2_X1 U284 ( .A(n194), .B(n319), .ZN(n271) );
  XNOR2_X1 U285 ( .A(n203), .B(n319), .ZN(n279) );
  XNOR2_X1 U286 ( .A(n319), .B(FCU_IF_ID_6_10[3]), .ZN(n170) );
  XNOR2_X1 U287 ( .A(FCU_EX_MEM_11_15[3]), .B(FCU_ID_EX_11_15[3]), .ZN(n250)
         );
  XNOR2_X1 U288 ( .A(FCU_ID_EX_6_10[3]), .B(FCU_EX_MEM_11_15[3]), .ZN(n221) );
  XNOR2_X1 U289 ( .A(n307), .B(FCU_IF_ID_6_10[0]), .ZN(n165) );
  XNOR2_X1 U290 ( .A(FCU_ID_EX_6_10[0]), .B(n307), .ZN(n213) );
  XNOR2_X1 U291 ( .A(n193), .B(n320), .ZN(n269) );
  XNOR2_X1 U292 ( .A(n204), .B(n320), .ZN(n277) );
  XNOR2_X1 U293 ( .A(n80), .B(n320), .ZN(n173) );
  XNOR2_X1 U294 ( .A(FCU_EX_MEM_11_15[4]), .B(FCU_ID_EX_6_10[4]), .ZN(n222) );
  XNOR2_X1 U295 ( .A(FCU_EX_MEM_16_20[1]), .B(FCU_ID_EX_11_15[1]), .ZN(n259)
         );
  XNOR2_X1 U296 ( .A(FCU_ID_EX_6_10[1]), .B(FCU_EX_MEM_16_20[1]), .ZN(n214) );
  INV_X1 U297 ( .A(n246), .ZN(n164) );
  OAI21_X1 U298 ( .B1(n208), .B2(n287), .A(s_stall_mem), .ZN(n205) );
  INV_X1 U299 ( .A(n227), .ZN(n226) );
  OAI21_X1 U300 ( .B1(n244), .B2(n243), .A(s_stall_mem), .ZN(n227) );
endmodule


module WriteBack_Stage_NBIT_DATA32 ( WB_OpA, WB_OpB, WB_sel, WB_reduce, 
        WB_BYTE_half, WB_SGN_usg, WB_out );
  input [31:0] WB_OpA;
  input [31:0] WB_OpB;
  output [31:0] WB_out;
  input WB_sel, WB_reduce, WB_BYTE_half, WB_SGN_usg;

  wire   [31:0] s_tmp;

  Mux_NBit_2x1_NBIT_IN32_80 WB_MUX ( .port0(WB_OpA), .port1(WB_OpB), .sel(
        WB_sel), .portY(s_tmp) );
  Sign_Reducer_NBIT_data32 WB_SGB ( .SR_data_in(s_tmp), .SR_reduce(WB_reduce), 
        .SR_BYTE_half(WB_BYTE_half), .SR_SGN_usg(WB_SGN_usg), .SR_data_out(
        WB_out) );
endmodule


module Memory_Stage_NBIT_DATA32_NBIT_ADDRESS32 ( ME_data_in, ME_address, 
        ME_clk, ME_rst, ME_enable, ME_reduce, ME_BYTE_half, ME_data_to_mem, 
        ME_address_to_mem, ME_data_from_mem, ME_data_rd_out );
  input [31:0] ME_data_in;
  input [31:0] ME_address;
  output [31:0] ME_data_to_mem;
  output [31:0] ME_address_to_mem;
  input [31:0] ME_data_from_mem;
  output [31:0] ME_data_rd_out;
  input ME_clk, ME_rst, ME_enable, ME_reduce, ME_BYTE_half;

  assign ME_address_to_mem[31] = ME_address[31];
  assign ME_address_to_mem[30] = ME_address[30];
  assign ME_address_to_mem[29] = ME_address[29];
  assign ME_address_to_mem[28] = ME_address[28];
  assign ME_address_to_mem[27] = ME_address[27];
  assign ME_address_to_mem[26] = ME_address[26];
  assign ME_address_to_mem[25] = ME_address[25];
  assign ME_address_to_mem[24] = ME_address[24];
  assign ME_address_to_mem[23] = ME_address[23];
  assign ME_address_to_mem[22] = ME_address[22];
  assign ME_address_to_mem[21] = ME_address[21];
  assign ME_address_to_mem[20] = ME_address[20];
  assign ME_address_to_mem[19] = ME_address[19];
  assign ME_address_to_mem[18] = ME_address[18];
  assign ME_address_to_mem[17] = ME_address[17];
  assign ME_address_to_mem[16] = ME_address[16];
  assign ME_address_to_mem[15] = ME_address[15];
  assign ME_address_to_mem[14] = ME_address[14];
  assign ME_address_to_mem[13] = ME_address[13];
  assign ME_address_to_mem[12] = ME_address[12];
  assign ME_address_to_mem[11] = ME_address[11];
  assign ME_address_to_mem[10] = ME_address[10];
  assign ME_address_to_mem[9] = ME_address[9];
  assign ME_address_to_mem[8] = ME_address[8];
  assign ME_address_to_mem[7] = ME_address[7];
  assign ME_address_to_mem[6] = ME_address[6];
  assign ME_address_to_mem[5] = ME_address[5];
  assign ME_address_to_mem[4] = ME_address[4];
  assign ME_address_to_mem[3] = ME_address[3];
  assign ME_address_to_mem[2] = ME_address[2];
  assign ME_address_to_mem[1] = ME_address[1];
  assign ME_address_to_mem[0] = ME_address[0];

  Data_Reducer_NBIT_DATA32 DR ( .DR_data_in(ME_data_in), .DR_reduce(ME_reduce), 
        .DR_BYTE_half(ME_BYTE_half), .DR_data_out(ME_data_to_mem) );
  NRegister_N32_33 REG_RD ( .clk(ME_clk), .reset(ME_rst), .data_in(
        ME_data_from_mem), .enable(ME_enable), .load(1'b1), .data_out(
        ME_data_rd_out) );
endmodule


module Execute_Stage_NBIT_DATA32_NBIT_BS_AMOUNT5 ( EX_clk, EX_reset, EX_enable, 
        EX_OpA, EX_OpB, EX_Opcode, EX_ShiftAmount, EX_sel_mux_out, EX_data_out, 
        EX_PSW );
  input [31:0] EX_OpA;
  input [31:0] EX_OpB;
  input [5:0] EX_Opcode;
  input [4:0] EX_ShiftAmount;
  input [1:0] EX_sel_mux_out;
  output [31:0] EX_data_out;
  output [4:0] EX_PSW;
  input EX_clk, EX_reset, EX_enable;
  wire   s_mul_enable, \s_mux_signals[1][0][31] , \s_mux_signals[1][0][30] ,
         \s_mux_signals[1][0][29] , \s_mux_signals[1][0][28] ,
         \s_mux_signals[1][0][27] , \s_mux_signals[1][0][26] ,
         \s_mux_signals[1][0][25] , \s_mux_signals[1][0][24] ,
         \s_mux_signals[1][0][23] , \s_mux_signals[1][0][22] ,
         \s_mux_signals[1][0][21] , \s_mux_signals[1][0][20] ,
         \s_mux_signals[1][0][19] , \s_mux_signals[1][0][18] ,
         \s_mux_signals[1][0][17] , \s_mux_signals[1][0][16] ,
         \s_mux_signals[1][0][15] , \s_mux_signals[1][0][14] ,
         \s_mux_signals[1][0][13] , \s_mux_signals[1][0][12] ,
         \s_mux_signals[1][0][11] , \s_mux_signals[1][0][10] ,
         \s_mux_signals[1][0][9] , \s_mux_signals[1][0][8] ,
         \s_mux_signals[1][0][7] , \s_mux_signals[1][0][6] ,
         \s_mux_signals[1][0][5] , \s_mux_signals[1][0][4] ,
         \s_mux_signals[1][0][3] , \s_mux_signals[1][0][2] ,
         \s_mux_signals[1][0][1] , \s_mux_signals[1][0][0] ,
         \s_mux_signals[1][1][31] , \s_mux_signals[1][1][30] ,
         \s_mux_signals[1][1][29] , \s_mux_signals[1][1][28] ,
         \s_mux_signals[1][1][27] , \s_mux_signals[1][1][26] ,
         \s_mux_signals[1][1][25] , \s_mux_signals[1][1][24] ,
         \s_mux_signals[1][1][23] , \s_mux_signals[1][1][22] ,
         \s_mux_signals[1][1][21] , \s_mux_signals[1][1][20] ,
         \s_mux_signals[1][1][19] , \s_mux_signals[1][1][18] ,
         \s_mux_signals[1][1][17] , \s_mux_signals[1][1][16] ,
         \s_mux_signals[1][1][15] , \s_mux_signals[1][1][14] ,
         \s_mux_signals[1][1][13] , \s_mux_signals[1][1][12] ,
         \s_mux_signals[1][1][11] , \s_mux_signals[1][1][10] ,
         \s_mux_signals[1][1][9] , \s_mux_signals[1][1][8] ,
         \s_mux_signals[1][1][7] , \s_mux_signals[1][1][6] ,
         \s_mux_signals[1][1][5] , \s_mux_signals[1][1][4] ,
         \s_mux_signals[1][1][3] , \s_mux_signals[1][1][2] ,
         \s_mux_signals[1][1][1] , \s_mux_signals[1][1][0] , n1, n3, n4, n5,
         n6, n7, n8, n9;
  wire   [31:0] s_OpA_Fei_Talu;
  wire   [31:0] s_OpB_Fei_Talu;
  wire   [31:0] s_OpA_Fei_Tmul;
  wire   [31:0] s_OpB_Fei_Tmul;
  wire   [31:0] s_outalu_Falu_Treg;
  wire   [4:0] s_flags_Falu_statusreg;
  wire   [63:0] s_product_Fmul_Thiloregs;
  wire   [31:0] s_product_Flo_Tmux;
  wire   [31:0] s_product_Fhi_Tmux;
  wire   [31:0] s_outalu_Falu_Tmux;

  Enable_Interface_NBIT_DATA32_0 EI_OpA_Alu ( .EI_datain({EX_OpA[31:2], n6, n7}), .EI_enable(n1), .EI_dataout(s_OpA_Fei_Talu) );
  Enable_Interface_NBIT_DATA32_3 EI_OpB_Alu ( .EI_datain({EX_OpB[31], n8, n5, 
        EX_OpB[28], n4, EX_OpB[26:0]}), .EI_enable(n1), .EI_dataout(
        s_OpB_Fei_Talu) );
  Enable_Interface_NBIT_DATA32_2 EI_OpA_Mul ( .EI_datain({n9, EX_OpA[30:0]}), 
        .EI_enable(s_mul_enable), .EI_dataout(s_OpA_Fei_Tmul) );
  Enable_Interface_NBIT_DATA32_1 EI_OpB_Mul ( .EI_datain(EX_OpB), .EI_enable(
        s_mul_enable), .EI_dataout(s_OpB_Fei_Tmul) );
  ALU_NBIT_ALU32_NBIT_BS_AMOUNT5 ALU_NBIT ( .ALU_OpA(s_OpA_Fei_Talu), 
        .ALU_OpB(s_OpB_Fei_Talu), .ALU_Opcode(EX_Opcode), .ALU_BS_amount(
        EX_ShiftAmount), .ALU_output(s_outalu_Falu_Treg), .ALU_flags(
        s_flags_Falu_statusreg) );
  Multiplier_NBIT_DATA32 MUL ( .MUL_OpA(s_OpA_Fei_Tmul), .MUL_OpB(
        s_OpB_Fei_Tmul), .MUL_SGN_usgn(EX_Opcode[1]), .MUL_product(
        s_product_Fmul_Thiloregs) );
  NRegister_N32_36 LO ( .clk(EX_clk), .reset(EX_reset), .data_in(
        s_product_Fmul_Thiloregs[31:0]), .enable(s_mul_enable), .load(1'b1), 
        .data_out(s_product_Flo_Tmux) );
  NRegister_N32_35 HI ( .clk(EX_clk), .reset(EX_reset), .data_in(
        s_product_Fmul_Thiloregs[63:32]), .enable(s_mul_enable), .load(1'b1), 
        .data_out(s_product_Fhi_Tmux) );
  NRegister_N32_34 ALU_reg ( .clk(EX_clk), .reset(EX_reset), .data_in(
        s_outalu_Falu_Treg), .enable(n1), .load(1'b1), .data_out(
        s_outalu_Falu_Tmux) );
  Mux_NBit_2x1_NBIT_IN32_83 MUX1 ( .port0(s_outalu_Falu_Tmux), .port1(
        s_product_Fhi_Tmux), .sel(EX_sel_mux_out[0]), .portY({
        \s_mux_signals[1][0][31] , \s_mux_signals[1][0][30] , 
        \s_mux_signals[1][0][29] , \s_mux_signals[1][0][28] , 
        \s_mux_signals[1][0][27] , \s_mux_signals[1][0][26] , 
        \s_mux_signals[1][0][25] , \s_mux_signals[1][0][24] , 
        \s_mux_signals[1][0][23] , \s_mux_signals[1][0][22] , 
        \s_mux_signals[1][0][21] , \s_mux_signals[1][0][20] , 
        \s_mux_signals[1][0][19] , \s_mux_signals[1][0][18] , 
        \s_mux_signals[1][0][17] , \s_mux_signals[1][0][16] , 
        \s_mux_signals[1][0][15] , \s_mux_signals[1][0][14] , 
        \s_mux_signals[1][0][13] , \s_mux_signals[1][0][12] , 
        \s_mux_signals[1][0][11] , \s_mux_signals[1][0][10] , 
        \s_mux_signals[1][0][9] , \s_mux_signals[1][0][8] , 
        \s_mux_signals[1][0][7] , \s_mux_signals[1][0][6] , 
        \s_mux_signals[1][0][5] , \s_mux_signals[1][0][4] , 
        \s_mux_signals[1][0][3] , \s_mux_signals[1][0][2] , 
        \s_mux_signals[1][0][1] , \s_mux_signals[1][0][0] }) );
  Mux_NBit_2x1_NBIT_IN32_82 MUX2 ( .port0(s_product_Flo_Tmux), .port1({1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sel(EX_sel_mux_out[0]), 
        .portY({\s_mux_signals[1][1][31] , \s_mux_signals[1][1][30] , 
        \s_mux_signals[1][1][29] , \s_mux_signals[1][1][28] , 
        \s_mux_signals[1][1][27] , \s_mux_signals[1][1][26] , 
        \s_mux_signals[1][1][25] , \s_mux_signals[1][1][24] , 
        \s_mux_signals[1][1][23] , \s_mux_signals[1][1][22] , 
        \s_mux_signals[1][1][21] , \s_mux_signals[1][1][20] , 
        \s_mux_signals[1][1][19] , \s_mux_signals[1][1][18] , 
        \s_mux_signals[1][1][17] , \s_mux_signals[1][1][16] , 
        \s_mux_signals[1][1][15] , \s_mux_signals[1][1][14] , 
        \s_mux_signals[1][1][13] , \s_mux_signals[1][1][12] , 
        \s_mux_signals[1][1][11] , \s_mux_signals[1][1][10] , 
        \s_mux_signals[1][1][9] , \s_mux_signals[1][1][8] , 
        \s_mux_signals[1][1][7] , \s_mux_signals[1][1][6] , 
        \s_mux_signals[1][1][5] , \s_mux_signals[1][1][4] , 
        \s_mux_signals[1][1][3] , \s_mux_signals[1][1][2] , 
        \s_mux_signals[1][1][1] , \s_mux_signals[1][1][0] }) );
  Mux_NBit_2x1_NBIT_IN32_81 MUX3 ( .port0({\s_mux_signals[1][0][31] , 
        \s_mux_signals[1][0][30] , \s_mux_signals[1][0][29] , 
        \s_mux_signals[1][0][28] , \s_mux_signals[1][0][27] , 
        \s_mux_signals[1][0][26] , \s_mux_signals[1][0][25] , 
        \s_mux_signals[1][0][24] , \s_mux_signals[1][0][23] , 
        \s_mux_signals[1][0][22] , \s_mux_signals[1][0][21] , 
        \s_mux_signals[1][0][20] , \s_mux_signals[1][0][19] , 
        \s_mux_signals[1][0][18] , \s_mux_signals[1][0][17] , 
        \s_mux_signals[1][0][16] , \s_mux_signals[1][0][15] , 
        \s_mux_signals[1][0][14] , \s_mux_signals[1][0][13] , 
        \s_mux_signals[1][0][12] , \s_mux_signals[1][0][11] , 
        \s_mux_signals[1][0][10] , \s_mux_signals[1][0][9] , 
        \s_mux_signals[1][0][8] , \s_mux_signals[1][0][7] , 
        \s_mux_signals[1][0][6] , \s_mux_signals[1][0][5] , 
        \s_mux_signals[1][0][4] , \s_mux_signals[1][0][3] , 
        \s_mux_signals[1][0][2] , \s_mux_signals[1][0][1] , 
        \s_mux_signals[1][0][0] }), .port1({\s_mux_signals[1][1][31] , 
        \s_mux_signals[1][1][30] , \s_mux_signals[1][1][29] , 
        \s_mux_signals[1][1][28] , \s_mux_signals[1][1][27] , 
        \s_mux_signals[1][1][26] , \s_mux_signals[1][1][25] , 
        \s_mux_signals[1][1][24] , \s_mux_signals[1][1][23] , 
        \s_mux_signals[1][1][22] , \s_mux_signals[1][1][21] , 
        \s_mux_signals[1][1][20] , \s_mux_signals[1][1][19] , 
        \s_mux_signals[1][1][18] , \s_mux_signals[1][1][17] , 
        \s_mux_signals[1][1][16] , \s_mux_signals[1][1][15] , 
        \s_mux_signals[1][1][14] , \s_mux_signals[1][1][13] , 
        \s_mux_signals[1][1][12] , \s_mux_signals[1][1][11] , 
        \s_mux_signals[1][1][10] , \s_mux_signals[1][1][9] , 
        \s_mux_signals[1][1][8] , \s_mux_signals[1][1][7] , 
        \s_mux_signals[1][1][6] , \s_mux_signals[1][1][5] , 
        \s_mux_signals[1][1][4] , \s_mux_signals[1][1][3] , 
        \s_mux_signals[1][1][2] , \s_mux_signals[1][1][1] , 
        \s_mux_signals[1][1][0] }), .sel(EX_sel_mux_out[1]), .portY(
        EX_data_out) );
  NRegister_N5_1 PSW ( .clk(EX_clk), .reset(EX_reset), .data_in(
        s_flags_Falu_statusreg), .enable(n1), .load(1'b1), .data_out(EX_PSW)
         );
  CLKBUF_X1 U3 ( .A(EX_OpB[27]), .Z(n4) );
  CLKBUF_X1 U4 ( .A(EX_OpB[29]), .Z(n5) );
  CLKBUF_X1 U5 ( .A(EX_OpA[1]), .Z(n6) );
  CLKBUF_X1 U6 ( .A(EX_OpA[0]), .Z(n7) );
  CLKBUF_X1 U7 ( .A(EX_OpB[30]), .Z(n8) );
  AOI21_X1 U8 ( .B1(EX_Opcode[5]), .B2(EX_Opcode[4]), .A(n3), .ZN(n1) );
  INV_X1 U9 ( .A(EX_enable), .ZN(n3) );
  AND3_X1 U10 ( .A1(EX_enable), .A2(EX_Opcode[4]), .A3(EX_Opcode[5]), .ZN(
        s_mul_enable) );
  CLKBUF_X1 U11 ( .A(EX_OpA[31]), .Z(n9) );
endmodule


module Mux_NBit_2x1_NBIT_IN5_3 ( port0, port1, sel, portY );
  input [4:0] port0;
  input [4:0] port1;
  output [4:0] portY;
  input sel;
  wire   N2, N3, N4, N6, n7, n8, n9, n10, n11, n12;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[4] = N6;

  INV_X1 U1 ( .A(n11), .ZN(N3) );
  INV_X1 U2 ( .A(n10), .ZN(N4) );
  AOI22_X1 U3 ( .A1(port0[2]), .A2(n8), .B1(port1[2]), .B2(sel), .ZN(n10) );
  AOI22_X1 U4 ( .A1(port0[1]), .A2(n8), .B1(port1[1]), .B2(sel), .ZN(n11) );
  AOI22_X1 U5 ( .A1(port0[0]), .A2(n8), .B1(port1[0]), .B2(sel), .ZN(n12) );
  AOI22_X1 U6 ( .A1(port0[4]), .A2(n8), .B1(port1[4]), .B2(sel), .ZN(n9) );
  INV_X1 U7 ( .A(sel), .ZN(n8) );
  INV_X1 U8 ( .A(n9), .ZN(N6) );
  INV_X1 U9 ( .A(n12), .ZN(N2) );
  INV_X1 U10 ( .A(n7), .ZN(portY[3]) );
  AOI22_X1 U11 ( .A1(port0[3]), .A2(n8), .B1(sel), .B2(port1[3]), .ZN(n7) );
endmodule


module Mux_NBit_2x1_NBIT_IN5_0 ( port0, port1, sel, portY );
  input [4:0] port0;
  input [4:0] port1;
  output [4:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, n7, n9, n10, n11, n12, n1, n2, n3;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;

  CLKBUF_X1 U1 ( .A(sel), .Z(n1) );
  CLKBUF_X1 U2 ( .A(sel), .Z(n2) );
  INV_X1 U3 ( .A(n11), .ZN(N3) );
  AOI22_X1 U4 ( .A1(port0[4]), .A2(n3), .B1(n2), .B2(port1[4]), .ZN(n7) );
  AOI22_X1 U5 ( .A1(port0[3]), .A2(n3), .B1(port1[3]), .B2(n1), .ZN(n9) );
  INV_X1 U6 ( .A(n12), .ZN(N2) );
  INV_X1 U7 ( .A(n9), .ZN(N5) );
  INV_X1 U8 ( .A(n7), .ZN(N6) );
  INV_X1 U9 ( .A(n10), .ZN(N4) );
  AOI22_X1 U10 ( .A1(port0[2]), .A2(n3), .B1(port1[2]), .B2(n1), .ZN(n10) );
  AOI22_X1 U11 ( .A1(port0[0]), .A2(n3), .B1(port1[0]), .B2(n1), .ZN(n12) );
  AOI22_X1 U12 ( .A1(port0[1]), .A2(n3), .B1(port1[1]), .B2(n1), .ZN(n11) );
  INV_X1 U13 ( .A(n2), .ZN(n3) );
endmodule


module Mux_NBit_2x1_NBIT_IN32_0 ( port0, port1, sel, portY );
  input [31:0] port0;
  input [31:0] port1;
  output [31:0] portY;
  input sel;
  wire   N2, N3, N4, N5, N6, N7, N8, N9, N10, N11, N12, N13, N14, N15, N16,
         N17, N18, N19, N20, N21, N22, N23, N24, N25, N26, N27, N28, N29, N30,
         N31, N32, N33, n34, n36, n37, n38, n39, n40, n41, n42, n43, n44, n45,
         n46, n47, n48, n49, n50, n51, n52, n53, n54, n55, n56, n57, n58, n59,
         n60, n61, n62, n63, n64, n65, n66, n1, n2, n3, n4, n5, n6, n7, n8, n9,
         n10, n11, n12, n13, n14, n15;
  assign portY[0] = N2;
  assign portY[1] = N3;
  assign portY[2] = N4;
  assign portY[3] = N5;
  assign portY[4] = N6;
  assign portY[5] = N7;
  assign portY[6] = N8;
  assign portY[7] = N9;
  assign portY[8] = N10;
  assign portY[9] = N11;
  assign portY[10] = N12;
  assign portY[11] = N13;
  assign portY[12] = N14;
  assign portY[13] = N15;
  assign portY[14] = N16;
  assign portY[15] = N17;
  assign portY[16] = N18;
  assign portY[17] = N19;
  assign portY[18] = N20;
  assign portY[19] = N21;
  assign portY[20] = N22;
  assign portY[21] = N23;
  assign portY[22] = N24;
  assign portY[23] = N25;
  assign portY[24] = N26;
  assign portY[25] = N27;
  assign portY[26] = N28;
  assign portY[27] = N29;
  assign portY[28] = N30;
  assign portY[29] = N31;
  assign portY[30] = N32;
  assign portY[31] = N33;

  CLKBUF_X1 U1 ( .A(n3), .Z(n14) );
  BUF_X1 U2 ( .A(n2), .Z(n12) );
  BUF_X1 U3 ( .A(n3), .Z(n15) );
  INV_X1 U4 ( .A(n15), .ZN(n5) );
  INV_X1 U5 ( .A(n15), .ZN(n4) );
  BUF_X1 U6 ( .A(n1), .Z(n8) );
  CLKBUF_X1 U7 ( .A(n1), .Z(n9) );
  BUF_X1 U8 ( .A(n2), .Z(n11) );
  CLKBUF_X1 U9 ( .A(n2), .Z(n10) );
  BUF_X1 U10 ( .A(n3), .Z(n13) );
  CLKBUF_X1 U11 ( .A(n1), .Z(n7) );
  BUF_X1 U12 ( .A(sel), .Z(n3) );
  CLKBUF_X1 U13 ( .A(sel), .Z(n1) );
  CLKBUF_X1 U14 ( .A(sel), .Z(n2) );
  INV_X1 U15 ( .A(n37), .ZN(N7) );
  AOI22_X1 U16 ( .A1(port0[5]), .A2(n6), .B1(port1[5]), .B2(n7), .ZN(n37) );
  INV_X1 U17 ( .A(n38), .ZN(N6) );
  AOI22_X1 U18 ( .A1(port0[4]), .A2(n6), .B1(port1[4]), .B2(n7), .ZN(n38) );
  INV_X1 U19 ( .A(n36), .ZN(N8) );
  AOI22_X1 U20 ( .A1(port0[6]), .A2(n6), .B1(port1[6]), .B2(n7), .ZN(n36) );
  INV_X1 U21 ( .A(n39), .ZN(N5) );
  AOI22_X1 U22 ( .A1(port0[3]), .A2(n6), .B1(port1[3]), .B2(n7), .ZN(n39) );
  INV_X1 U23 ( .A(n42), .ZN(N32) );
  AOI22_X1 U24 ( .A1(port0[30]), .A2(n6), .B1(port1[30]), .B2(n8), .ZN(n42) );
  INV_X1 U25 ( .A(n34), .ZN(N9) );
  AOI22_X1 U26 ( .A1(port0[7]), .A2(n6), .B1(n14), .B2(port1[7]), .ZN(n34) );
  INV_X1 U27 ( .A(n40), .ZN(N4) );
  AOI22_X1 U28 ( .A1(port0[2]), .A2(n6), .B1(port1[2]), .B2(n8), .ZN(n40) );
  INV_X1 U29 ( .A(n47), .ZN(N28) );
  AOI22_X1 U30 ( .A1(port0[26]), .A2(n5), .B1(port1[26]), .B2(n9), .ZN(n47) );
  INV_X1 U31 ( .A(n51), .ZN(N24) );
  AOI22_X1 U32 ( .A1(port0[22]), .A2(n5), .B1(port1[22]), .B2(n10), .ZN(n51)
         );
  INV_X1 U33 ( .A(n52), .ZN(N23) );
  AOI22_X1 U34 ( .A1(port0[21]), .A2(n5), .B1(port1[21]), .B2(n10), .ZN(n52)
         );
  INV_X1 U35 ( .A(n43), .ZN(N31) );
  AOI22_X1 U36 ( .A1(port0[29]), .A2(n5), .B1(port1[29]), .B2(n11), .ZN(n43)
         );
  INV_X1 U37 ( .A(n60), .ZN(N16) );
  AOI22_X1 U38 ( .A1(port0[14]), .A2(n4), .B1(port1[14]), .B2(n13), .ZN(n60)
         );
  INV_X1 U39 ( .A(n50), .ZN(N25) );
  AOI22_X1 U40 ( .A1(port0[23]), .A2(n5), .B1(port1[23]), .B2(n10), .ZN(n50)
         );
  INV_X1 U41 ( .A(n44), .ZN(N30) );
  AOI22_X1 U42 ( .A1(port0[28]), .A2(n5), .B1(port1[28]), .B2(n8), .ZN(n44) );
  INV_X1 U43 ( .A(n53), .ZN(N22) );
  AOI22_X1 U44 ( .A1(port0[20]), .A2(n5), .B1(port1[20]), .B2(n11), .ZN(n53)
         );
  INV_X1 U45 ( .A(n59), .ZN(N17) );
  AOI22_X1 U46 ( .A1(port0[15]), .A2(n4), .B1(port1[15]), .B2(n12), .ZN(n59)
         );
  INV_X1 U47 ( .A(n61), .ZN(N15) );
  AOI22_X1 U48 ( .A1(port0[13]), .A2(n4), .B1(port1[13]), .B2(n13), .ZN(n61)
         );
  INV_X1 U49 ( .A(n54), .ZN(N21) );
  AOI22_X1 U50 ( .A1(port0[19]), .A2(n5), .B1(port1[19]), .B2(n11), .ZN(n54)
         );
  INV_X1 U51 ( .A(n66), .ZN(N10) );
  AOI22_X1 U52 ( .A1(port0[8]), .A2(n4), .B1(port1[8]), .B2(n14), .ZN(n66) );
  INV_X1 U53 ( .A(n62), .ZN(N14) );
  AOI22_X1 U54 ( .A1(port0[12]), .A2(n4), .B1(port1[12]), .B2(n13), .ZN(n62)
         );
  INV_X1 U55 ( .A(n64), .ZN(N12) );
  AOI22_X1 U56 ( .A1(port0[10]), .A2(n4), .B1(port1[10]), .B2(n14), .ZN(n64)
         );
  INV_X1 U57 ( .A(n63), .ZN(N13) );
  AOI22_X1 U58 ( .A1(port0[11]), .A2(n4), .B1(port1[11]), .B2(n13), .ZN(n63)
         );
  INV_X1 U59 ( .A(n46), .ZN(N29) );
  AOI22_X1 U60 ( .A1(port0[27]), .A2(n5), .B1(port1[27]), .B2(n9), .ZN(n46) );
  INV_X1 U61 ( .A(n65), .ZN(N11) );
  AOI22_X1 U62 ( .A1(port0[9]), .A2(n4), .B1(port1[9]), .B2(n14), .ZN(n65) );
  INV_X1 U63 ( .A(n49), .ZN(N26) );
  AOI22_X1 U64 ( .A1(port0[24]), .A2(n5), .B1(port1[24]), .B2(n10), .ZN(n49)
         );
  INV_X1 U65 ( .A(n45), .ZN(N3) );
  AOI22_X1 U66 ( .A1(port0[1]), .A2(n5), .B1(port1[1]), .B2(n9), .ZN(n45) );
  INV_X1 U67 ( .A(n55), .ZN(N20) );
  AOI22_X1 U68 ( .A1(port0[18]), .A2(n4), .B1(port1[18]), .B2(n11), .ZN(n55)
         );
  INV_X1 U69 ( .A(n58), .ZN(N18) );
  AOI22_X1 U70 ( .A1(port0[16]), .A2(n4), .B1(port1[16]), .B2(n12), .ZN(n58)
         );
  INV_X1 U71 ( .A(n57), .ZN(N19) );
  AOI22_X1 U72 ( .A1(port0[17]), .A2(n4), .B1(port1[17]), .B2(n12), .ZN(n57)
         );
  INV_X1 U73 ( .A(n48), .ZN(N27) );
  AOI22_X1 U74 ( .A1(port0[25]), .A2(n5), .B1(port1[25]), .B2(n9), .ZN(n48) );
  INV_X1 U75 ( .A(n56), .ZN(N2) );
  AOI22_X1 U76 ( .A1(port0[0]), .A2(n4), .B1(port1[0]), .B2(n12), .ZN(n56) );
  INV_X1 U77 ( .A(n41), .ZN(N33) );
  AOI22_X1 U78 ( .A1(port0[31]), .A2(n6), .B1(port1[31]), .B2(n8), .ZN(n41) );
  INV_X1 U79 ( .A(n15), .ZN(n6) );
endmodule


module Decode_NBIT_PC32_NBIT_IR32_NBIT_ADDR5_NBIT_DATA32 ( DE_clk, DE_reset, 
        DE_enable, DE_stall, DE_IR, DE_PC, DE_NPC, DE_rd1, DE_rd2, DE_wr, 
        DE_data_fex, DE_sel_data_forward, DE_data_Fwb, DE_signext, 
        DE_JMP_branch, DE_jmp_or_branch, DE_save_PC, DE_branch_taken, 
        DE_new_PC, DE_imm_address, DE_RegA, DE_RegB, DE_RegI );
  input [31:0] DE_IR;
  input [31:0] DE_PC;
  input [31:0] DE_NPC;
  input [31:0] DE_data_fex;
  input [1:0] DE_sel_data_forward;
  input [31:0] DE_data_Fwb;
  input [1:0] DE_signext;
  input [1:0] DE_JMP_branch;
  output [31:0] DE_new_PC;
  output [31:0] DE_imm_address;
  output [31:0] DE_RegA;
  output [31:0] DE_RegB;
  output [31:0] DE_RegI;
  input DE_clk, DE_reset, DE_enable, DE_stall, DE_rd1, DE_rd2, DE_wr,
         DE_jmp_or_branch, DE_save_PC;
  output DE_branch_taken;
  wire   s_enable1, s_enable2, s_wr_de, s_wr_ex, s_wr_mem, s_notRd2,
         s_iszero_Fcmp_Tcond, s_prev_instr_branch_taken, s_isnt_jmp_or_branch,
         n3, n2, n4;
  wire   [4:0] s_wr_addr_type;
  wire   [4:0] s_fmux_tr1;
  wire   [4:0] s_ex;
  wire   [4:0] s_mem;
  wire   [4:0] s_wb;
  wire   [31:0] s_data_Frf_TregA;
  wire   [31:0] s_data_Frf_TregB;
  wire   [31:0] s_fwd_tmp;
  wire   [31:0] s_fwd_fmux_tcmp;

  Reg1Bit_7 R1_enable ( .clk(DE_clk), .reset(n4), .data_in(DE_stall), .enable(
        DE_enable), .load(1'b1), .data_out(s_enable1) );
  Reg1Bit_6 R2_enable ( .clk(DE_clk), .reset(n4), .data_in(s_enable1), 
        .enable(DE_enable), .load(1'b1), .data_out(s_enable2) );
  Reg1Bit_5 R3_enable ( .clk(DE_clk), .reset(n4), .data_in(s_enable2), 
        .enable(DE_enable), .load(1'b1) );
  Reg1Bit_4 R1_wr ( .clk(DE_clk), .reset(n4), .data_in(DE_wr), .enable(
        DE_stall), .load(1'b1), .data_out(s_wr_de) );
  Reg1Bit_3 R2_wr ( .clk(DE_clk), .reset(n4), .data_in(s_wr_de), .enable(
        s_enable1), .load(1'b1), .data_out(s_wr_ex) );
  Reg1Bit_2 R3_wr ( .clk(DE_clk), .reset(n4), .data_in(s_wr_ex), .enable(
        s_enable2), .load(1'b1), .data_out(s_wr_mem) );
  Mux_NBit_2x1_NBIT_IN5_2 TypeWr_MUX ( .port0(DE_IR[15:11]), .port1(
        DE_IR[20:16]), .sel(s_notRd2), .portY(s_wr_addr_type) );
  Mux_NBit_2x1_NBIT_IN5_1 Write_MUX ( .port0(s_wr_addr_type), .port1({1'b1, 
        1'b1, 1'b1, 1'b1, 1'b1}), .sel(DE_save_PC), .portY(s_fmux_tr1) );
  NRegister_N5_0 R1 ( .clk(DE_clk), .reset(n4), .data_in(s_fmux_tr1), .enable(
        DE_stall), .load(1'b1), .data_out(s_ex) );
  NRegister_N5_3 R2 ( .clk(DE_clk), .reset(n4), .data_in(s_ex), .enable(
        s_enable1), .load(1'b1), .data_out(s_mem) );
  NRegister_N5_2 R3 ( .clk(DE_clk), .reset(n4), .data_in(s_mem), .enable(
        s_enable2), .load(1'b1), .data_out(s_wb) );
  Register_File_NBIT_ADDR5_NBIT_DATA32 RF ( .RF_clk(DE_clk), .RF_reset(n4), 
        .RF_enable(DE_enable), .RF_RD1(DE_rd1), .RF_RD2(DE_rd2), .RF_WR(
        s_wr_mem), .RF_AddrRd1(DE_IR[25:21]), .RF_AddrRd2(DE_IR[20:16]), 
        .RF_AddrWr(s_wb), .RF_data_in(DE_data_Fwb), .RF_out1(s_data_Frf_TregA), 
        .RF_out2(s_data_Frf_TregB) );
  Sign_Extender_NBIT_DATA32 SE ( .SE_I_J(DE_signext[1]), .SE_S_U(DE_signext[0]), .SE_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, DE_IR[25:0]}), .SE_out(
        DE_imm_address) );
  Mux_NBit_2x1_NBIT_IN32_85 FWD_MUX1 ( .port0({s_data_Frf_TregA[31:1], n2}), 
        .port1(DE_data_fex), .sel(DE_sel_data_forward[0]), .portY(s_fwd_tmp)
         );
  Mux_NBit_2x1_NBIT_IN32_84 FWD_MUX2 ( .port0(s_fwd_tmp), .port1(DE_data_Fwb), 
        .sel(DE_sel_data_forward[1]), .portY(s_fwd_fmux_tcmp) );
  NRegister_N32_39 RegA ( .clk(DE_clk), .reset(n4), .data_in({
        s_data_Frf_TregA[31:1], n2}), .enable(DE_enable), .load(1'b1), 
        .data_out(DE_RegA) );
  NRegister_N32_38 RegB ( .clk(DE_clk), .reset(n4), .data_in(s_data_Frf_TregB), 
        .enable(DE_enable), .load(1'b1), .data_out(DE_RegB) );
  NRegister_N32_37 RegI ( .clk(DE_clk), .reset(n4), .data_in(DE_imm_address), 
        .enable(DE_enable), .load(1'b1), .data_out(DE_RegI) );
  NComparatorWithEnable_NBIT32_1 Cmp ( .A(s_fwd_fmux_tcmp), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Enable(DE_enable), 
        .ComparatorBit(s_iszero_Fcmp_Tcond) );
  Jmp_Branch_Manager_N32 JBM ( .JBM_iszero(s_iszero_Fcmp_Tcond), .JBM_Reg(
        s_data_Frf_TregA), .JBM_Imm(DE_imm_address), .JBM_NPC(DE_NPC), 
        .JBM_JMP_branch(DE_JMP_branch), .JBM_transparent_mode(
        s_isnt_jmp_or_branch), .JBM_Upd_PC(DE_new_PC), .JBM_taken(
        DE_branch_taken) );
  Reg1Bit_1 Branch_taken_reg ( .clk(DE_clk), .reset(n4), .data_in(
        DE_branch_taken), .enable(DE_stall), .load(1'b1), .data_out(
        s_prev_instr_branch_taken) );
  CLKBUF_X1 U3 ( .A(s_data_Frf_TregA[0]), .Z(n2) );
  BUF_X1 U4 ( .A(DE_reset), .Z(n4) );
  NAND2_X1 U5 ( .A1(DE_jmp_or_branch), .A2(n3), .ZN(s_isnt_jmp_or_branch) );
  INV_X1 U6 ( .A(s_prev_instr_branch_taken), .ZN(n3) );
  INV_X1 U7 ( .A(DE_rd2), .ZN(s_notRd2) );
endmodule


module Reg1Bit_23 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n2, net106835, n6, n7, n4, n5;

  DFFR_X1 data_out_reg ( .D(n2), .CK(clk), .RN(n5), .Q(data_out), .QN(
        net106835) );
  OAI22_X1 U3 ( .A1(net106835), .A2(n6), .B1(n7), .B2(n4), .ZN(n2) );
  INV_X1 U4 ( .A(n7), .ZN(n6) );
  NAND2_X1 U5 ( .A1(load), .A2(enable), .ZN(n7) );
  INV_X1 U6 ( .A(data_in), .ZN(n4) );
  INV_X1 U7 ( .A(reset), .ZN(n5) );
endmodule


module NRegister_N32_117 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108226, net108227, net108228, net108229, net108230,
         net108231, net108232, net108233, net108234, net108235, net108236,
         net108237, net108238, net108239, net108240, net108241, net108242,
         net108243, net108244, net108245, net108246, net108247, net108248,
         net108249, net108250, net108251, net108252, net108253, net108254,
         net108255, net108256, net108257, n68, n69, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n46), .Q(data_out[31]), 
        .QN(net108257) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n44), .Q(data_out[30]), 
        .QN(net108256) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n44), .Q(data_out[29]), 
        .QN(net108255) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n44), .Q(data_out[28]), 
        .QN(net108254) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n44), .Q(data_out[27]), 
        .QN(net108253) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n44), .Q(data_out[26]), 
        .QN(net108252) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n44), .Q(data_out[25]), 
        .QN(net108251) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n46), .Q(data_out[24]), 
        .QN(net108250) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n44), .Q(data_out[23]), 
        .QN(net108249) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n45), .Q(data_out[22]), 
        .QN(net108248) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n45), .Q(data_out[21]), 
        .QN(net108247) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n45), .Q(data_out[20]), 
        .QN(net108246) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n45), .Q(data_out[19]), 
        .QN(net108245) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n45), .Q(data_out[18]), 
        .QN(net108244) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n45), .Q(data_out[17]), 
        .QN(net108243) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n45), .Q(data_out[16]), 
        .QN(net108242) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n44), .Q(data_out[15]), 
        .QN(net108241) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n46), .Q(data_out[14]), 
        .QN(net108240) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n44), .Q(data_out[13]), 
        .QN(net108239) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108238) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108237) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n44), .Q(data_out[10]), 
        .QN(net108236) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n44), .Q(data_out[9]), 
        .QN(net108235) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n44), .Q(data_out[8]), 
        .QN(net108234) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108233) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n45), .Q(data_out[6]), 
        .QN(net108232) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n45), .Q(data_out[5]), 
        .QN(net108231) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n46), .Q(data_out[4]), 
        .QN(net108230) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n46), .Q(data_out[3]), 
        .QN(net108229) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n46), .Q(data_out[2]), 
        .QN(net108228) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n46), .Q(data_out[1]), 
        .QN(net108227) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n46), .Q(data_out[0]), 
        .QN(net108226) );
  BUF_X1 U3 ( .A(n47), .Z(n45) );
  BUF_X1 U4 ( .A(n47), .Z(n44) );
  BUF_X1 U5 ( .A(n47), .Z(n46) );
  INV_X1 U6 ( .A(n43), .ZN(n35) );
  INV_X1 U7 ( .A(reset), .ZN(n47) );
  BUF_X1 U8 ( .A(n68), .Z(n39) );
  BUF_X1 U9 ( .A(n68), .Z(n40) );
  BUF_X1 U10 ( .A(n68), .Z(n42) );
  BUF_X1 U11 ( .A(n68), .Z(n37) );
  BUF_X1 U12 ( .A(n68), .Z(n38) );
  BUF_X1 U13 ( .A(n68), .Z(n41) );
  BUF_X1 U14 ( .A(n68), .Z(n43) );
  OAI22_X1 U15 ( .A1(n37), .A2(n74), .B1(net108255), .B2(n36), .ZN(n5) );
  INV_X1 U16 ( .A(data_in[29]), .ZN(n74) );
  OAI22_X1 U17 ( .A1(n37), .A2(n73), .B1(net108254), .B2(n36), .ZN(n6) );
  INV_X1 U18 ( .A(data_in[28]), .ZN(n73) );
  OAI22_X1 U19 ( .A1(n37), .A2(n72), .B1(net108253), .B2(n36), .ZN(n7) );
  INV_X1 U20 ( .A(data_in[27]), .ZN(n72) );
  OAI22_X1 U21 ( .A1(n37), .A2(n71), .B1(net108252), .B2(n36), .ZN(n8) );
  INV_X1 U22 ( .A(data_in[26]), .ZN(n71) );
  OAI22_X1 U23 ( .A1(n91), .A2(n41), .B1(net108257), .B2(n35), .ZN(n2) );
  INV_X1 U24 ( .A(data_in[31]), .ZN(n91) );
  OAI22_X1 U25 ( .A1(n38), .A2(n75), .B1(net108256), .B2(n36), .ZN(n4) );
  INV_X1 U26 ( .A(data_in[30]), .ZN(n75) );
  OAI22_X1 U27 ( .A1(n37), .A2(n69), .B1(net108251), .B2(n36), .ZN(n9) );
  INV_X1 U28 ( .A(data_in[25]), .ZN(n69) );
  OAI22_X1 U29 ( .A1(n38), .A2(n76), .B1(net108226), .B2(n36), .ZN(n34) );
  INV_X1 U30 ( .A(data_in[0]), .ZN(n76) );
  OAI22_X1 U31 ( .A1(n38), .A2(n77), .B1(net108227), .B2(n36), .ZN(n33) );
  INV_X1 U32 ( .A(data_in[1]), .ZN(n77) );
  OAI22_X1 U33 ( .A1(n43), .A2(n101), .B1(net108250), .B2(n35), .ZN(n10) );
  INV_X1 U34 ( .A(data_in[24]), .ZN(n101) );
  OAI22_X1 U35 ( .A1(n43), .A2(n100), .B1(net108249), .B2(n35), .ZN(n11) );
  INV_X1 U36 ( .A(data_in[23]), .ZN(n100) );
  OAI22_X1 U37 ( .A1(n42), .A2(n99), .B1(net108248), .B2(n35), .ZN(n12) );
  INV_X1 U38 ( .A(data_in[22]), .ZN(n99) );
  OAI22_X1 U39 ( .A1(n42), .A2(n98), .B1(net108247), .B2(n35), .ZN(n13) );
  INV_X1 U40 ( .A(data_in[21]), .ZN(n98) );
  OAI22_X1 U41 ( .A1(n42), .A2(n97), .B1(net108246), .B2(n35), .ZN(n14) );
  INV_X1 U42 ( .A(data_in[20]), .ZN(n97) );
  OAI22_X1 U43 ( .A1(n42), .A2(n96), .B1(net108245), .B2(n35), .ZN(n15) );
  INV_X1 U44 ( .A(data_in[19]), .ZN(n96) );
  OAI22_X1 U45 ( .A1(n42), .A2(n95), .B1(net108244), .B2(n35), .ZN(n16) );
  INV_X1 U46 ( .A(data_in[18]), .ZN(n95) );
  OAI22_X1 U47 ( .A1(n40), .A2(n88), .B1(net108238), .B2(n35), .ZN(n22) );
  INV_X1 U48 ( .A(data_in[12]), .ZN(n88) );
  OAI22_X1 U49 ( .A1(n40), .A2(n89), .B1(net108239), .B2(n36), .ZN(n21) );
  INV_X1 U50 ( .A(data_in[13]), .ZN(n89) );
  OAI22_X1 U51 ( .A1(n41), .A2(n90), .B1(net108240), .B2(n35), .ZN(n20) );
  INV_X1 U52 ( .A(data_in[14]), .ZN(n90) );
  OAI22_X1 U53 ( .A1(n41), .A2(n94), .B1(net108243), .B2(n35), .ZN(n17) );
  INV_X1 U54 ( .A(data_in[17]), .ZN(n94) );
  OAI22_X1 U55 ( .A1(n41), .A2(n93), .B1(net108242), .B2(n35), .ZN(n18) );
  INV_X1 U56 ( .A(data_in[16]), .ZN(n93) );
  OAI22_X1 U57 ( .A1(n41), .A2(n92), .B1(net108241), .B2(n35), .ZN(n19) );
  INV_X1 U58 ( .A(data_in[15]), .ZN(n92) );
  OAI22_X1 U59 ( .A1(n39), .A2(n84), .B1(net108234), .B2(n35), .ZN(n26) );
  INV_X1 U60 ( .A(data_in[8]), .ZN(n84) );
  OAI22_X1 U61 ( .A1(n40), .A2(n85), .B1(net108235), .B2(n36), .ZN(n25) );
  INV_X1 U62 ( .A(data_in[9]), .ZN(n85) );
  OAI22_X1 U63 ( .A1(n40), .A2(n86), .B1(net108236), .B2(n35), .ZN(n24) );
  INV_X1 U64 ( .A(data_in[10]), .ZN(n86) );
  OAI22_X1 U65 ( .A1(n40), .A2(n87), .B1(net108237), .B2(n36), .ZN(n23) );
  INV_X1 U66 ( .A(data_in[11]), .ZN(n87) );
  OAI22_X1 U67 ( .A1(n38), .A2(n78), .B1(net108228), .B2(n35), .ZN(n32) );
  INV_X1 U68 ( .A(data_in[2]), .ZN(n78) );
  OAI22_X1 U69 ( .A1(n38), .A2(n79), .B1(net108229), .B2(n36), .ZN(n31) );
  INV_X1 U70 ( .A(data_in[3]), .ZN(n79) );
  OAI22_X1 U71 ( .A1(n39), .A2(n80), .B1(net108230), .B2(n36), .ZN(n30) );
  INV_X1 U72 ( .A(data_in[4]), .ZN(n80) );
  OAI22_X1 U73 ( .A1(n39), .A2(n81), .B1(net108231), .B2(n36), .ZN(n29) );
  INV_X1 U74 ( .A(data_in[5]), .ZN(n81) );
  OAI22_X1 U75 ( .A1(n39), .A2(n82), .B1(net108232), .B2(n36), .ZN(n28) );
  INV_X1 U76 ( .A(data_in[6]), .ZN(n82) );
  OAI22_X1 U77 ( .A1(n39), .A2(n83), .B1(net108233), .B2(n36), .ZN(n27) );
  INV_X1 U78 ( .A(data_in[7]), .ZN(n83) );
  NAND2_X1 U79 ( .A1(load), .A2(enable), .ZN(n68) );
  INV_X1 U80 ( .A(n43), .ZN(n36) );
endmodule


module NRegister_N32_118 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n2, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16, n17,
         n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31,
         n32, n33, n34, net108194, net108195, net108196, net108197, net108198,
         net108199, net108200, net108201, net108202, net108203, net108204,
         net108205, net108206, net108207, net108208, net108209, net108210,
         net108211, net108212, net108213, net108214, net108215, net108216,
         net108217, net108218, net108219, net108220, net108221, net108222,
         net108223, net108224, net108225, n68, n69, n71, n72, n73, n74, n75,
         n76, n77, n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89,
         n90, n91, n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47;

  DFFR_X1 \data_out_reg[31]  ( .D(n2), .CK(clk), .RN(n46), .Q(data_out[31]), 
        .QN(net108225) );
  DFFR_X1 \data_out_reg[30]  ( .D(n4), .CK(clk), .RN(n46), .Q(data_out[30]), 
        .QN(net108224) );
  DFFR_X1 \data_out_reg[29]  ( .D(n5), .CK(clk), .RN(n46), .Q(data_out[29]), 
        .QN(net108223) );
  DFFR_X1 \data_out_reg[28]  ( .D(n6), .CK(clk), .RN(n44), .Q(data_out[28]), 
        .QN(net108222) );
  DFFR_X1 \data_out_reg[27]  ( .D(n7), .CK(clk), .RN(n46), .Q(data_out[27]), 
        .QN(net108221) );
  DFFR_X1 \data_out_reg[26]  ( .D(n8), .CK(clk), .RN(n44), .Q(data_out[26]), 
        .QN(net108220) );
  DFFR_X1 \data_out_reg[25]  ( .D(n9), .CK(clk), .RN(n44), .Q(data_out[25]), 
        .QN(net108219) );
  DFFR_X1 \data_out_reg[24]  ( .D(n10), .CK(clk), .RN(n44), .Q(data_out[24]), 
        .QN(net108218) );
  DFFR_X1 \data_out_reg[23]  ( .D(n11), .CK(clk), .RN(n46), .Q(data_out[23]), 
        .QN(net108217) );
  DFFR_X1 \data_out_reg[22]  ( .D(n12), .CK(clk), .RN(n44), .Q(data_out[22]), 
        .QN(net108216) );
  DFFR_X1 \data_out_reg[21]  ( .D(n13), .CK(clk), .RN(n44), .Q(data_out[21]), 
        .QN(net108215) );
  DFFR_X1 \data_out_reg[20]  ( .D(n14), .CK(clk), .RN(n44), .Q(data_out[20]), 
        .QN(net108214) );
  DFFR_X1 \data_out_reg[19]  ( .D(n15), .CK(clk), .RN(n44), .Q(data_out[19]), 
        .QN(net108213) );
  DFFR_X1 \data_out_reg[18]  ( .D(n16), .CK(clk), .RN(n44), .Q(data_out[18]), 
        .QN(net108212) );
  DFFR_X1 \data_out_reg[17]  ( .D(n17), .CK(clk), .RN(n44), .Q(data_out[17]), 
        .QN(net108211) );
  DFFR_X1 \data_out_reg[16]  ( .D(n18), .CK(clk), .RN(n44), .Q(data_out[16]), 
        .QN(net108210) );
  DFFR_X1 \data_out_reg[15]  ( .D(n19), .CK(clk), .RN(n44), .Q(data_out[15]), 
        .QN(net108209) );
  DFFR_X1 \data_out_reg[14]  ( .D(n20), .CK(clk), .RN(n45), .Q(data_out[14]), 
        .QN(net108208) );
  DFFR_X1 \data_out_reg[13]  ( .D(n21), .CK(clk), .RN(n45), .Q(data_out[13]), 
        .QN(net108207) );
  DFFR_X1 \data_out_reg[12]  ( .D(n22), .CK(clk), .RN(n45), .Q(data_out[12]), 
        .QN(net108206) );
  DFFR_X1 \data_out_reg[11]  ( .D(n23), .CK(clk), .RN(n45), .Q(data_out[11]), 
        .QN(net108205) );
  DFFR_X1 \data_out_reg[10]  ( .D(n24), .CK(clk), .RN(n45), .Q(data_out[10]), 
        .QN(net108204) );
  DFFR_X1 \data_out_reg[9]  ( .D(n25), .CK(clk), .RN(n45), .Q(data_out[9]), 
        .QN(net108203) );
  DFFR_X1 \data_out_reg[8]  ( .D(n26), .CK(clk), .RN(n45), .Q(data_out[8]), 
        .QN(net108202) );
  DFFR_X1 \data_out_reg[7]  ( .D(n27), .CK(clk), .RN(n45), .Q(data_out[7]), 
        .QN(net108201) );
  DFFR_X1 \data_out_reg[6]  ( .D(n28), .CK(clk), .RN(n45), .Q(data_out[6]), 
        .QN(net108200) );
  DFFR_X1 \data_out_reg[5]  ( .D(n29), .CK(clk), .RN(n45), .Q(data_out[5]), 
        .QN(net108199) );
  DFFR_X1 \data_out_reg[4]  ( .D(n30), .CK(clk), .RN(n45), .Q(data_out[4]), 
        .QN(net108198) );
  DFFR_X1 \data_out_reg[3]  ( .D(n31), .CK(clk), .RN(n45), .Q(data_out[3]), 
        .QN(net108197) );
  DFFR_X1 \data_out_reg[2]  ( .D(n32), .CK(clk), .RN(n46), .Q(data_out[2]), 
        .QN(net108196) );
  DFFR_X1 \data_out_reg[1]  ( .D(n33), .CK(clk), .RN(n46), .Q(data_out[1]), 
        .QN(net108195) );
  DFFR_X1 \data_out_reg[0]  ( .D(n34), .CK(clk), .RN(n46), .Q(data_out[0]), 
        .QN(net108194) );
  BUF_X1 U3 ( .A(n47), .Z(n45) );
  BUF_X1 U4 ( .A(n47), .Z(n44) );
  BUF_X1 U5 ( .A(n47), .Z(n46) );
  INV_X1 U6 ( .A(n43), .ZN(n36) );
  INV_X1 U7 ( .A(n43), .ZN(n35) );
  INV_X1 U8 ( .A(reset), .ZN(n47) );
  BUF_X1 U9 ( .A(n68), .Z(n39) );
  BUF_X1 U10 ( .A(n68), .Z(n40) );
  BUF_X1 U11 ( .A(n68), .Z(n42) );
  BUF_X1 U12 ( .A(n68), .Z(n37) );
  BUF_X1 U13 ( .A(n68), .Z(n38) );
  BUF_X1 U14 ( .A(n68), .Z(n41) );
  BUF_X1 U15 ( .A(n68), .Z(n43) );
  NAND2_X1 U16 ( .A1(load), .A2(enable), .ZN(n68) );
  OAI22_X1 U17 ( .A1(n38), .A2(n76), .B1(net108194), .B2(n36), .ZN(n34) );
  INV_X1 U18 ( .A(data_in[0]), .ZN(n76) );
  OAI22_X1 U19 ( .A1(n38), .A2(n77), .B1(net108195), .B2(n35), .ZN(n33) );
  INV_X1 U20 ( .A(data_in[1]), .ZN(n77) );
  OAI22_X1 U21 ( .A1(n37), .A2(n69), .B1(net108219), .B2(n36), .ZN(n9) );
  INV_X1 U22 ( .A(data_in[25]), .ZN(n69) );
  OAI22_X1 U23 ( .A1(n37), .A2(n71), .B1(net108220), .B2(n35), .ZN(n8) );
  INV_X1 U24 ( .A(data_in[26]), .ZN(n71) );
  OAI22_X1 U25 ( .A1(n37), .A2(n72), .B1(net108221), .B2(n36), .ZN(n7) );
  INV_X1 U26 ( .A(data_in[27]), .ZN(n72) );
  OAI22_X1 U27 ( .A1(n37), .A2(n73), .B1(net108222), .B2(n35), .ZN(n6) );
  INV_X1 U28 ( .A(data_in[28]), .ZN(n73) );
  OAI22_X1 U29 ( .A1(n37), .A2(n74), .B1(net108223), .B2(n36), .ZN(n5) );
  INV_X1 U30 ( .A(data_in[29]), .ZN(n74) );
  OAI22_X1 U31 ( .A1(n38), .A2(n75), .B1(net108224), .B2(n35), .ZN(n4) );
  INV_X1 U32 ( .A(data_in[30]), .ZN(n75) );
  OAI22_X1 U33 ( .A1(n38), .A2(n78), .B1(net108196), .B2(n36), .ZN(n32) );
  INV_X1 U34 ( .A(data_in[2]), .ZN(n78) );
  OAI22_X1 U35 ( .A1(n38), .A2(n79), .B1(net108197), .B2(n36), .ZN(n31) );
  INV_X1 U36 ( .A(data_in[3]), .ZN(n79) );
  OAI22_X1 U37 ( .A1(n39), .A2(n80), .B1(net108198), .B2(n36), .ZN(n30) );
  INV_X1 U38 ( .A(data_in[4]), .ZN(n80) );
  OAI22_X1 U39 ( .A1(n39), .A2(n81), .B1(net108199), .B2(n36), .ZN(n29) );
  INV_X1 U40 ( .A(data_in[5]), .ZN(n81) );
  OAI22_X1 U41 ( .A1(n39), .A2(n82), .B1(net108200), .B2(n36), .ZN(n28) );
  INV_X1 U42 ( .A(data_in[6]), .ZN(n82) );
  OAI22_X1 U43 ( .A1(n39), .A2(n83), .B1(net108201), .B2(n36), .ZN(n27) );
  INV_X1 U44 ( .A(data_in[7]), .ZN(n83) );
  OAI22_X1 U45 ( .A1(n39), .A2(n84), .B1(net108202), .B2(n36), .ZN(n26) );
  INV_X1 U46 ( .A(data_in[8]), .ZN(n84) );
  OAI22_X1 U47 ( .A1(n40), .A2(n85), .B1(net108203), .B2(n36), .ZN(n25) );
  INV_X1 U48 ( .A(data_in[9]), .ZN(n85) );
  OAI22_X1 U49 ( .A1(n40), .A2(n86), .B1(net108204), .B2(n36), .ZN(n24) );
  INV_X1 U50 ( .A(data_in[10]), .ZN(n86) );
  OAI22_X1 U51 ( .A1(n40), .A2(n87), .B1(net108205), .B2(n36), .ZN(n23) );
  INV_X1 U52 ( .A(data_in[11]), .ZN(n87) );
  OAI22_X1 U53 ( .A1(n40), .A2(n88), .B1(net108206), .B2(n36), .ZN(n22) );
  INV_X1 U54 ( .A(data_in[12]), .ZN(n88) );
  OAI22_X1 U55 ( .A1(n40), .A2(n89), .B1(net108207), .B2(n36), .ZN(n21) );
  INV_X1 U56 ( .A(data_in[13]), .ZN(n89) );
  OAI22_X1 U57 ( .A1(n41), .A2(n90), .B1(net108208), .B2(n35), .ZN(n20) );
  INV_X1 U58 ( .A(data_in[14]), .ZN(n90) );
  OAI22_X1 U59 ( .A1(n41), .A2(n92), .B1(net108209), .B2(n35), .ZN(n19) );
  INV_X1 U60 ( .A(data_in[15]), .ZN(n92) );
  OAI22_X1 U61 ( .A1(n41), .A2(n93), .B1(net108210), .B2(n35), .ZN(n18) );
  INV_X1 U62 ( .A(data_in[16]), .ZN(n93) );
  OAI22_X1 U63 ( .A1(n41), .A2(n94), .B1(net108211), .B2(n35), .ZN(n17) );
  INV_X1 U64 ( .A(data_in[17]), .ZN(n94) );
  OAI22_X1 U65 ( .A1(n42), .A2(n95), .B1(net108212), .B2(n35), .ZN(n16) );
  INV_X1 U66 ( .A(data_in[18]), .ZN(n95) );
  OAI22_X1 U67 ( .A1(n42), .A2(n96), .B1(net108213), .B2(n35), .ZN(n15) );
  INV_X1 U68 ( .A(data_in[19]), .ZN(n96) );
  OAI22_X1 U69 ( .A1(n42), .A2(n97), .B1(net108214), .B2(n35), .ZN(n14) );
  INV_X1 U70 ( .A(data_in[20]), .ZN(n97) );
  OAI22_X1 U71 ( .A1(n42), .A2(n98), .B1(net108215), .B2(n35), .ZN(n13) );
  INV_X1 U72 ( .A(data_in[21]), .ZN(n98) );
  OAI22_X1 U73 ( .A1(n42), .A2(n99), .B1(net108216), .B2(n35), .ZN(n12) );
  INV_X1 U74 ( .A(data_in[22]), .ZN(n99) );
  OAI22_X1 U75 ( .A1(n43), .A2(n100), .B1(net108217), .B2(n35), .ZN(n11) );
  INV_X1 U76 ( .A(data_in[23]), .ZN(n100) );
  OAI22_X1 U77 ( .A1(n43), .A2(n101), .B1(net108218), .B2(n35), .ZN(n10) );
  INV_X1 U78 ( .A(data_in[24]), .ZN(n101) );
  OAI22_X1 U79 ( .A1(n41), .A2(n91), .B1(net108225), .B2(n35), .ZN(n2) );
  INV_X1 U80 ( .A(data_in[31]), .ZN(n91) );
endmodule


module Fetch_NBIT_PC32_NBIT_IR32 ( FE_clk, FE_rst, FE_enable, FE_PC_enable, 
        FE_PC_clear, FE_IR_enable, FE_IR_clear, FE_btb_target_prediction, 
        FE_btb_prediction, FE_branch_taken, FE_next_instr_is_branch, 
        FE_next_instr_is_jump, FE_new_PC_from_DE, FE_IR_in, FE_restore_BTB, 
        FE_IR_out, FE_PC, FE_NPC );
  input [31:0] FE_btb_target_prediction;
  input [31:0] FE_new_PC_from_DE;
  input [31:0] FE_IR_in;
  output [31:0] FE_IR_out;
  output [31:0] FE_PC;
  output [31:0] FE_NPC;
  input FE_clk, FE_rst, FE_enable, FE_PC_enable, FE_PC_clear, FE_IR_enable,
         FE_IR_clear, FE_btb_prediction, FE_branch_taken,
         FE_next_instr_is_branch, FE_next_instr_is_jump;
  output FE_restore_BTB;
  wire   s_pc_rst, s_pc_enable, s_ir_rst, s_ir_enable, s_inc_sel,
         s_btb_prediction, s_jmp, n3, n5, n6, n7;
  wire   [31:0] s_tmp;
  wire   [31:0] s_sum_Fcla_Tnpcreg;
  wire   [31:0] s_restored_pc;
  wire   [31:0] s_target_Fbtbmux_Tnpcmux;
  wire   [31:0] s_tmp_pc;

  NRegister_N32_42 PC ( .clk(FE_clk), .reset(s_pc_rst), .data_in(FE_NPC), 
        .enable(s_pc_enable), .load(1'b1), .data_out(FE_PC) );
  NRegister_N32_41 IR ( .clk(FE_clk), .reset(s_ir_rst), .data_in(FE_IR_in), 
        .enable(s_ir_enable), .load(1'b1), .data_out(FE_IR_out) );
  Mux_NBit_2x1_NBIT_IN32_89 MUXN_INC ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .port1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b1, 1'b0, 
        1'b0}), .sel(s_inc_sel), .portY(s_tmp) );
  PropagateCarryLookahead_N32_0 ADDPC ( .A(FE_PC), .B(s_tmp), .Cin(1'b0), 
        .Sum(s_sum_Fcla_Tnpcreg) );
  NRegister_N32_40 Restore_PC ( .clk(FE_clk), .reset(s_pc_rst), .data_in(
        s_sum_Fcla_Tnpcreg), .enable(s_pc_enable), .load(1'b1), .data_out(
        s_restored_pc) );
  Mux_NBit_2x1_NBIT_IN32_88 MUXBTB ( .port0(s_sum_Fcla_Tnpcreg), .port1(
        FE_btb_target_prediction), .sel(FE_btb_prediction), .portY(
        s_target_Fbtbmux_Tnpcmux) );
  Reg1Bit_8 BTB_prediction_reg ( .clk(FE_clk), .reset(s_pc_rst), .data_in(
        FE_btb_prediction), .enable(s_pc_enable), .load(1'b1), .data_out(
        s_btb_prediction) );
  Mux_NBit_2x1_NBIT_IN32_87 MUXNPC ( .port0(s_target_Fbtbmux_Tnpcmux), .port1(
        FE_new_PC_from_DE), .sel(s_jmp), .portY(s_tmp_pc) );
  Mux_NBit_2x1_NBIT_IN32_86 MUX_restore ( .port0(s_tmp_pc), .port1(
        s_restored_pc), .sel(FE_restore_BTB), .portY(FE_NPC) );
  AND3_X2 U3 ( .A1(FE_next_instr_is_jump), .A2(n3), .A3(FE_branch_taken), .ZN(
        s_jmp) );
  NOR2_X1 U4 ( .A1(FE_rst), .A2(n7), .ZN(s_inc_sel) );
  AND2_X1 U5 ( .A1(n6), .A2(FE_PC_enable), .ZN(s_pc_enable) );
  OR2_X1 U6 ( .A1(FE_PC_clear), .A2(FE_rst), .ZN(s_pc_rst) );
  OR2_X1 U7 ( .A1(FE_IR_clear), .A2(FE_rst), .ZN(s_ir_rst) );
  NOR3_X1 U8 ( .A1(n3), .A2(FE_branch_taken), .A3(n5), .ZN(FE_restore_BTB) );
  INV_X1 U9 ( .A(FE_next_instr_is_jump), .ZN(n5) );
  AND2_X1 U10 ( .A1(FE_IR_enable), .A2(n6), .ZN(s_ir_enable) );
  NAND2_X1 U11 ( .A1(s_btb_prediction), .A2(FE_next_instr_is_branch), .ZN(n3)
         );
  INV_X1 U12 ( .A(n7), .ZN(n6) );
  INV_X1 U13 ( .A(FE_enable), .ZN(n7) );
endmodule


module BTB_N_ENTRY32_NBIT_ENTRY32_NBIT_TARGET32_NBIT_PREDICTION3 ( BTB_clk, 
        BTB_rst, BTB_enable, BTB_restore, BTB_PC_From_IF, BTB_PC_From_DE, 
        BTB_target_From_DE, BTB_is_branch, BTB_branch_taken, 
        BTB_target_prediction, BTB_prediction );
  input [31:0] BTB_PC_From_IF;
  input [31:0] BTB_PC_From_DE;
  input [31:0] BTB_target_From_DE;
  output [31:0] BTB_target_prediction;
  input BTB_clk, BTB_rst, BTB_enable, BTB_restore, BTB_is_branch,
         BTB_branch_taken;
  output BTB_prediction;
  wire   \s_entries_Freg_Tcmp[0][31] , \s_entries_Freg_Tcmp[0][30] ,
         \s_entries_Freg_Tcmp[0][29] , \s_entries_Freg_Tcmp[0][28] ,
         \s_entries_Freg_Tcmp[0][27] , \s_entries_Freg_Tcmp[0][26] ,
         \s_entries_Freg_Tcmp[0][25] , \s_entries_Freg_Tcmp[0][24] ,
         \s_entries_Freg_Tcmp[0][23] , \s_entries_Freg_Tcmp[0][22] ,
         \s_entries_Freg_Tcmp[0][21] , \s_entries_Freg_Tcmp[0][20] ,
         \s_entries_Freg_Tcmp[0][19] , \s_entries_Freg_Tcmp[0][18] ,
         \s_entries_Freg_Tcmp[0][17] , \s_entries_Freg_Tcmp[0][16] ,
         \s_entries_Freg_Tcmp[0][15] , \s_entries_Freg_Tcmp[0][14] ,
         \s_entries_Freg_Tcmp[0][13] , \s_entries_Freg_Tcmp[0][12] ,
         \s_entries_Freg_Tcmp[0][11] , \s_entries_Freg_Tcmp[0][10] ,
         \s_entries_Freg_Tcmp[0][9] , \s_entries_Freg_Tcmp[0][8] ,
         \s_entries_Freg_Tcmp[0][7] , \s_entries_Freg_Tcmp[0][6] ,
         \s_entries_Freg_Tcmp[0][5] , \s_entries_Freg_Tcmp[0][4] ,
         \s_entries_Freg_Tcmp[0][3] , \s_entries_Freg_Tcmp[0][2] ,
         \s_entries_Freg_Tcmp[0][1] , \s_entries_Freg_Tcmp[0][0] ,
         \s_entries_Freg_Tcmp[1][31] , \s_entries_Freg_Tcmp[1][30] ,
         \s_entries_Freg_Tcmp[1][29] , \s_entries_Freg_Tcmp[1][28] ,
         \s_entries_Freg_Tcmp[1][27] , \s_entries_Freg_Tcmp[1][26] ,
         \s_entries_Freg_Tcmp[1][25] , \s_entries_Freg_Tcmp[1][24] ,
         \s_entries_Freg_Tcmp[1][23] , \s_entries_Freg_Tcmp[1][22] ,
         \s_entries_Freg_Tcmp[1][21] , \s_entries_Freg_Tcmp[1][20] ,
         \s_entries_Freg_Tcmp[1][19] , \s_entries_Freg_Tcmp[1][18] ,
         \s_entries_Freg_Tcmp[1][17] , \s_entries_Freg_Tcmp[1][16] ,
         \s_entries_Freg_Tcmp[1][15] , \s_entries_Freg_Tcmp[1][14] ,
         \s_entries_Freg_Tcmp[1][13] , \s_entries_Freg_Tcmp[1][12] ,
         \s_entries_Freg_Tcmp[1][11] , \s_entries_Freg_Tcmp[1][10] ,
         \s_entries_Freg_Tcmp[1][9] , \s_entries_Freg_Tcmp[1][8] ,
         \s_entries_Freg_Tcmp[1][7] , \s_entries_Freg_Tcmp[1][6] ,
         \s_entries_Freg_Tcmp[1][5] , \s_entries_Freg_Tcmp[1][4] ,
         \s_entries_Freg_Tcmp[1][3] , \s_entries_Freg_Tcmp[1][2] ,
         \s_entries_Freg_Tcmp[1][1] , \s_entries_Freg_Tcmp[1][0] ,
         \s_entries_Freg_Tcmp[2][31] , \s_entries_Freg_Tcmp[2][30] ,
         \s_entries_Freg_Tcmp[2][29] , \s_entries_Freg_Tcmp[2][28] ,
         \s_entries_Freg_Tcmp[2][27] , \s_entries_Freg_Tcmp[2][26] ,
         \s_entries_Freg_Tcmp[2][25] , \s_entries_Freg_Tcmp[2][24] ,
         \s_entries_Freg_Tcmp[2][23] , \s_entries_Freg_Tcmp[2][22] ,
         \s_entries_Freg_Tcmp[2][21] , \s_entries_Freg_Tcmp[2][20] ,
         \s_entries_Freg_Tcmp[2][19] , \s_entries_Freg_Tcmp[2][18] ,
         \s_entries_Freg_Tcmp[2][17] , \s_entries_Freg_Tcmp[2][16] ,
         \s_entries_Freg_Tcmp[2][15] , \s_entries_Freg_Tcmp[2][14] ,
         \s_entries_Freg_Tcmp[2][13] , \s_entries_Freg_Tcmp[2][12] ,
         \s_entries_Freg_Tcmp[2][11] , \s_entries_Freg_Tcmp[2][10] ,
         \s_entries_Freg_Tcmp[2][9] , \s_entries_Freg_Tcmp[2][8] ,
         \s_entries_Freg_Tcmp[2][7] , \s_entries_Freg_Tcmp[2][6] ,
         \s_entries_Freg_Tcmp[2][5] , \s_entries_Freg_Tcmp[2][4] ,
         \s_entries_Freg_Tcmp[2][3] , \s_entries_Freg_Tcmp[2][2] ,
         \s_entries_Freg_Tcmp[2][1] , \s_entries_Freg_Tcmp[2][0] ,
         \s_entries_Freg_Tcmp[3][31] , \s_entries_Freg_Tcmp[3][30] ,
         \s_entries_Freg_Tcmp[3][29] , \s_entries_Freg_Tcmp[3][28] ,
         \s_entries_Freg_Tcmp[3][27] , \s_entries_Freg_Tcmp[3][26] ,
         \s_entries_Freg_Tcmp[3][25] , \s_entries_Freg_Tcmp[3][24] ,
         \s_entries_Freg_Tcmp[3][23] , \s_entries_Freg_Tcmp[3][22] ,
         \s_entries_Freg_Tcmp[3][21] , \s_entries_Freg_Tcmp[3][20] ,
         \s_entries_Freg_Tcmp[3][19] , \s_entries_Freg_Tcmp[3][18] ,
         \s_entries_Freg_Tcmp[3][17] , \s_entries_Freg_Tcmp[3][16] ,
         \s_entries_Freg_Tcmp[3][15] , \s_entries_Freg_Tcmp[3][14] ,
         \s_entries_Freg_Tcmp[3][13] , \s_entries_Freg_Tcmp[3][12] ,
         \s_entries_Freg_Tcmp[3][11] , \s_entries_Freg_Tcmp[3][10] ,
         \s_entries_Freg_Tcmp[3][9] , \s_entries_Freg_Tcmp[3][8] ,
         \s_entries_Freg_Tcmp[3][7] , \s_entries_Freg_Tcmp[3][6] ,
         \s_entries_Freg_Tcmp[3][5] , \s_entries_Freg_Tcmp[3][4] ,
         \s_entries_Freg_Tcmp[3][3] , \s_entries_Freg_Tcmp[3][2] ,
         \s_entries_Freg_Tcmp[3][1] , \s_entries_Freg_Tcmp[3][0] ,
         \s_entries_Freg_Tcmp[4][31] , \s_entries_Freg_Tcmp[4][30] ,
         \s_entries_Freg_Tcmp[4][29] , \s_entries_Freg_Tcmp[4][28] ,
         \s_entries_Freg_Tcmp[4][27] , \s_entries_Freg_Tcmp[4][26] ,
         \s_entries_Freg_Tcmp[4][25] , \s_entries_Freg_Tcmp[4][24] ,
         \s_entries_Freg_Tcmp[4][23] , \s_entries_Freg_Tcmp[4][22] ,
         \s_entries_Freg_Tcmp[4][21] , \s_entries_Freg_Tcmp[4][20] ,
         \s_entries_Freg_Tcmp[4][19] , \s_entries_Freg_Tcmp[4][18] ,
         \s_entries_Freg_Tcmp[4][17] , \s_entries_Freg_Tcmp[4][16] ,
         \s_entries_Freg_Tcmp[4][15] , \s_entries_Freg_Tcmp[4][14] ,
         \s_entries_Freg_Tcmp[4][13] , \s_entries_Freg_Tcmp[4][12] ,
         \s_entries_Freg_Tcmp[4][11] , \s_entries_Freg_Tcmp[4][10] ,
         \s_entries_Freg_Tcmp[4][9] , \s_entries_Freg_Tcmp[4][8] ,
         \s_entries_Freg_Tcmp[4][7] , \s_entries_Freg_Tcmp[4][6] ,
         \s_entries_Freg_Tcmp[4][5] , \s_entries_Freg_Tcmp[4][4] ,
         \s_entries_Freg_Tcmp[4][3] , \s_entries_Freg_Tcmp[4][2] ,
         \s_entries_Freg_Tcmp[4][1] , \s_entries_Freg_Tcmp[4][0] ,
         \s_entries_Freg_Tcmp[5][31] , \s_entries_Freg_Tcmp[5][30] ,
         \s_entries_Freg_Tcmp[5][29] , \s_entries_Freg_Tcmp[5][28] ,
         \s_entries_Freg_Tcmp[5][27] , \s_entries_Freg_Tcmp[5][26] ,
         \s_entries_Freg_Tcmp[5][25] , \s_entries_Freg_Tcmp[5][24] ,
         \s_entries_Freg_Tcmp[5][23] , \s_entries_Freg_Tcmp[5][22] ,
         \s_entries_Freg_Tcmp[5][21] , \s_entries_Freg_Tcmp[5][20] ,
         \s_entries_Freg_Tcmp[5][19] , \s_entries_Freg_Tcmp[5][18] ,
         \s_entries_Freg_Tcmp[5][17] , \s_entries_Freg_Tcmp[5][16] ,
         \s_entries_Freg_Tcmp[5][15] , \s_entries_Freg_Tcmp[5][14] ,
         \s_entries_Freg_Tcmp[5][13] , \s_entries_Freg_Tcmp[5][12] ,
         \s_entries_Freg_Tcmp[5][11] , \s_entries_Freg_Tcmp[5][10] ,
         \s_entries_Freg_Tcmp[5][9] , \s_entries_Freg_Tcmp[5][8] ,
         \s_entries_Freg_Tcmp[5][7] , \s_entries_Freg_Tcmp[5][6] ,
         \s_entries_Freg_Tcmp[5][5] , \s_entries_Freg_Tcmp[5][4] ,
         \s_entries_Freg_Tcmp[5][3] , \s_entries_Freg_Tcmp[5][2] ,
         \s_entries_Freg_Tcmp[5][1] , \s_entries_Freg_Tcmp[5][0] ,
         \s_entries_Freg_Tcmp[6][31] , \s_entries_Freg_Tcmp[6][30] ,
         \s_entries_Freg_Tcmp[6][29] , \s_entries_Freg_Tcmp[6][28] ,
         \s_entries_Freg_Tcmp[6][27] , \s_entries_Freg_Tcmp[6][26] ,
         \s_entries_Freg_Tcmp[6][25] , \s_entries_Freg_Tcmp[6][24] ,
         \s_entries_Freg_Tcmp[6][23] , \s_entries_Freg_Tcmp[6][22] ,
         \s_entries_Freg_Tcmp[6][21] , \s_entries_Freg_Tcmp[6][20] ,
         \s_entries_Freg_Tcmp[6][19] , \s_entries_Freg_Tcmp[6][18] ,
         \s_entries_Freg_Tcmp[6][17] , \s_entries_Freg_Tcmp[6][16] ,
         \s_entries_Freg_Tcmp[6][15] , \s_entries_Freg_Tcmp[6][14] ,
         \s_entries_Freg_Tcmp[6][13] , \s_entries_Freg_Tcmp[6][12] ,
         \s_entries_Freg_Tcmp[6][11] , \s_entries_Freg_Tcmp[6][10] ,
         \s_entries_Freg_Tcmp[6][9] , \s_entries_Freg_Tcmp[6][8] ,
         \s_entries_Freg_Tcmp[6][7] , \s_entries_Freg_Tcmp[6][6] ,
         \s_entries_Freg_Tcmp[6][5] , \s_entries_Freg_Tcmp[6][4] ,
         \s_entries_Freg_Tcmp[6][3] , \s_entries_Freg_Tcmp[6][2] ,
         \s_entries_Freg_Tcmp[6][1] , \s_entries_Freg_Tcmp[6][0] ,
         \s_entries_Freg_Tcmp[7][31] , \s_entries_Freg_Tcmp[7][30] ,
         \s_entries_Freg_Tcmp[7][29] , \s_entries_Freg_Tcmp[7][28] ,
         \s_entries_Freg_Tcmp[7][27] , \s_entries_Freg_Tcmp[7][26] ,
         \s_entries_Freg_Tcmp[7][25] , \s_entries_Freg_Tcmp[7][24] ,
         \s_entries_Freg_Tcmp[7][23] , \s_entries_Freg_Tcmp[7][22] ,
         \s_entries_Freg_Tcmp[7][21] , \s_entries_Freg_Tcmp[7][20] ,
         \s_entries_Freg_Tcmp[7][19] , \s_entries_Freg_Tcmp[7][18] ,
         \s_entries_Freg_Tcmp[7][17] , \s_entries_Freg_Tcmp[7][16] ,
         \s_entries_Freg_Tcmp[7][15] , \s_entries_Freg_Tcmp[7][14] ,
         \s_entries_Freg_Tcmp[7][13] , \s_entries_Freg_Tcmp[7][12] ,
         \s_entries_Freg_Tcmp[7][11] , \s_entries_Freg_Tcmp[7][10] ,
         \s_entries_Freg_Tcmp[7][9] , \s_entries_Freg_Tcmp[7][8] ,
         \s_entries_Freg_Tcmp[7][7] , \s_entries_Freg_Tcmp[7][6] ,
         \s_entries_Freg_Tcmp[7][5] , \s_entries_Freg_Tcmp[7][4] ,
         \s_entries_Freg_Tcmp[7][3] , \s_entries_Freg_Tcmp[7][2] ,
         \s_entries_Freg_Tcmp[7][1] , \s_entries_Freg_Tcmp[7][0] ,
         \s_entries_Freg_Tcmp[8][31] , \s_entries_Freg_Tcmp[8][30] ,
         \s_entries_Freg_Tcmp[8][29] , \s_entries_Freg_Tcmp[8][28] ,
         \s_entries_Freg_Tcmp[8][27] , \s_entries_Freg_Tcmp[8][26] ,
         \s_entries_Freg_Tcmp[8][25] , \s_entries_Freg_Tcmp[8][24] ,
         \s_entries_Freg_Tcmp[8][23] , \s_entries_Freg_Tcmp[8][22] ,
         \s_entries_Freg_Tcmp[8][21] , \s_entries_Freg_Tcmp[8][20] ,
         \s_entries_Freg_Tcmp[8][19] , \s_entries_Freg_Tcmp[8][18] ,
         \s_entries_Freg_Tcmp[8][17] , \s_entries_Freg_Tcmp[8][16] ,
         \s_entries_Freg_Tcmp[8][15] , \s_entries_Freg_Tcmp[8][14] ,
         \s_entries_Freg_Tcmp[8][13] , \s_entries_Freg_Tcmp[8][12] ,
         \s_entries_Freg_Tcmp[8][11] , \s_entries_Freg_Tcmp[8][10] ,
         \s_entries_Freg_Tcmp[8][9] , \s_entries_Freg_Tcmp[8][8] ,
         \s_entries_Freg_Tcmp[8][7] , \s_entries_Freg_Tcmp[8][6] ,
         \s_entries_Freg_Tcmp[8][5] , \s_entries_Freg_Tcmp[8][4] ,
         \s_entries_Freg_Tcmp[8][3] , \s_entries_Freg_Tcmp[8][2] ,
         \s_entries_Freg_Tcmp[8][1] , \s_entries_Freg_Tcmp[8][0] ,
         \s_entries_Freg_Tcmp[9][31] , \s_entries_Freg_Tcmp[9][30] ,
         \s_entries_Freg_Tcmp[9][29] , \s_entries_Freg_Tcmp[9][28] ,
         \s_entries_Freg_Tcmp[9][27] , \s_entries_Freg_Tcmp[9][26] ,
         \s_entries_Freg_Tcmp[9][25] , \s_entries_Freg_Tcmp[9][24] ,
         \s_entries_Freg_Tcmp[9][23] , \s_entries_Freg_Tcmp[9][22] ,
         \s_entries_Freg_Tcmp[9][21] , \s_entries_Freg_Tcmp[9][20] ,
         \s_entries_Freg_Tcmp[9][19] , \s_entries_Freg_Tcmp[9][18] ,
         \s_entries_Freg_Tcmp[9][17] , \s_entries_Freg_Tcmp[9][16] ,
         \s_entries_Freg_Tcmp[9][15] , \s_entries_Freg_Tcmp[9][14] ,
         \s_entries_Freg_Tcmp[9][13] , \s_entries_Freg_Tcmp[9][12] ,
         \s_entries_Freg_Tcmp[9][11] , \s_entries_Freg_Tcmp[9][10] ,
         \s_entries_Freg_Tcmp[9][9] , \s_entries_Freg_Tcmp[9][8] ,
         \s_entries_Freg_Tcmp[9][7] , \s_entries_Freg_Tcmp[9][6] ,
         \s_entries_Freg_Tcmp[9][5] , \s_entries_Freg_Tcmp[9][4] ,
         \s_entries_Freg_Tcmp[9][3] , \s_entries_Freg_Tcmp[9][2] ,
         \s_entries_Freg_Tcmp[9][1] , \s_entries_Freg_Tcmp[9][0] ,
         \s_entries_Freg_Tcmp[10][31] , \s_entries_Freg_Tcmp[10][30] ,
         \s_entries_Freg_Tcmp[10][29] , \s_entries_Freg_Tcmp[10][28] ,
         \s_entries_Freg_Tcmp[10][27] , \s_entries_Freg_Tcmp[10][26] ,
         \s_entries_Freg_Tcmp[10][25] , \s_entries_Freg_Tcmp[10][24] ,
         \s_entries_Freg_Tcmp[10][23] , \s_entries_Freg_Tcmp[10][22] ,
         \s_entries_Freg_Tcmp[10][21] , \s_entries_Freg_Tcmp[10][20] ,
         \s_entries_Freg_Tcmp[10][19] , \s_entries_Freg_Tcmp[10][18] ,
         \s_entries_Freg_Tcmp[10][17] , \s_entries_Freg_Tcmp[10][16] ,
         \s_entries_Freg_Tcmp[10][15] , \s_entries_Freg_Tcmp[10][14] ,
         \s_entries_Freg_Tcmp[10][13] , \s_entries_Freg_Tcmp[10][12] ,
         \s_entries_Freg_Tcmp[10][11] , \s_entries_Freg_Tcmp[10][10] ,
         \s_entries_Freg_Tcmp[10][9] , \s_entries_Freg_Tcmp[10][8] ,
         \s_entries_Freg_Tcmp[10][7] , \s_entries_Freg_Tcmp[10][6] ,
         \s_entries_Freg_Tcmp[10][5] , \s_entries_Freg_Tcmp[10][4] ,
         \s_entries_Freg_Tcmp[10][3] , \s_entries_Freg_Tcmp[10][2] ,
         \s_entries_Freg_Tcmp[10][1] , \s_entries_Freg_Tcmp[10][0] ,
         \s_entries_Freg_Tcmp[11][31] , \s_entries_Freg_Tcmp[11][30] ,
         \s_entries_Freg_Tcmp[11][29] , \s_entries_Freg_Tcmp[11][28] ,
         \s_entries_Freg_Tcmp[11][27] , \s_entries_Freg_Tcmp[11][26] ,
         \s_entries_Freg_Tcmp[11][25] , \s_entries_Freg_Tcmp[11][24] ,
         \s_entries_Freg_Tcmp[11][23] , \s_entries_Freg_Tcmp[11][22] ,
         \s_entries_Freg_Tcmp[11][21] , \s_entries_Freg_Tcmp[11][20] ,
         \s_entries_Freg_Tcmp[11][19] , \s_entries_Freg_Tcmp[11][18] ,
         \s_entries_Freg_Tcmp[11][17] , \s_entries_Freg_Tcmp[11][16] ,
         \s_entries_Freg_Tcmp[11][15] , \s_entries_Freg_Tcmp[11][14] ,
         \s_entries_Freg_Tcmp[11][13] , \s_entries_Freg_Tcmp[11][12] ,
         \s_entries_Freg_Tcmp[11][11] , \s_entries_Freg_Tcmp[11][10] ,
         \s_entries_Freg_Tcmp[11][9] , \s_entries_Freg_Tcmp[11][8] ,
         \s_entries_Freg_Tcmp[11][7] , \s_entries_Freg_Tcmp[11][6] ,
         \s_entries_Freg_Tcmp[11][5] , \s_entries_Freg_Tcmp[11][4] ,
         \s_entries_Freg_Tcmp[11][3] , \s_entries_Freg_Tcmp[11][2] ,
         \s_entries_Freg_Tcmp[11][1] , \s_entries_Freg_Tcmp[11][0] ,
         \s_entries_Freg_Tcmp[12][31] , \s_entries_Freg_Tcmp[12][30] ,
         \s_entries_Freg_Tcmp[12][29] , \s_entries_Freg_Tcmp[12][28] ,
         \s_entries_Freg_Tcmp[12][27] , \s_entries_Freg_Tcmp[12][26] ,
         \s_entries_Freg_Tcmp[12][25] , \s_entries_Freg_Tcmp[12][24] ,
         \s_entries_Freg_Tcmp[12][23] , \s_entries_Freg_Tcmp[12][22] ,
         \s_entries_Freg_Tcmp[12][21] , \s_entries_Freg_Tcmp[12][20] ,
         \s_entries_Freg_Tcmp[12][19] , \s_entries_Freg_Tcmp[12][18] ,
         \s_entries_Freg_Tcmp[12][17] , \s_entries_Freg_Tcmp[12][16] ,
         \s_entries_Freg_Tcmp[12][15] , \s_entries_Freg_Tcmp[12][14] ,
         \s_entries_Freg_Tcmp[12][13] , \s_entries_Freg_Tcmp[12][12] ,
         \s_entries_Freg_Tcmp[12][11] , \s_entries_Freg_Tcmp[12][10] ,
         \s_entries_Freg_Tcmp[12][9] , \s_entries_Freg_Tcmp[12][8] ,
         \s_entries_Freg_Tcmp[12][7] , \s_entries_Freg_Tcmp[12][6] ,
         \s_entries_Freg_Tcmp[12][5] , \s_entries_Freg_Tcmp[12][4] ,
         \s_entries_Freg_Tcmp[12][3] , \s_entries_Freg_Tcmp[12][2] ,
         \s_entries_Freg_Tcmp[12][1] , \s_entries_Freg_Tcmp[12][0] ,
         \s_entries_Freg_Tcmp[13][31] , \s_entries_Freg_Tcmp[13][30] ,
         \s_entries_Freg_Tcmp[13][29] , \s_entries_Freg_Tcmp[13][28] ,
         \s_entries_Freg_Tcmp[13][27] , \s_entries_Freg_Tcmp[13][26] ,
         \s_entries_Freg_Tcmp[13][25] , \s_entries_Freg_Tcmp[13][24] ,
         \s_entries_Freg_Tcmp[13][23] , \s_entries_Freg_Tcmp[13][22] ,
         \s_entries_Freg_Tcmp[13][21] , \s_entries_Freg_Tcmp[13][20] ,
         \s_entries_Freg_Tcmp[13][19] , \s_entries_Freg_Tcmp[13][18] ,
         \s_entries_Freg_Tcmp[13][17] , \s_entries_Freg_Tcmp[13][16] ,
         \s_entries_Freg_Tcmp[13][15] , \s_entries_Freg_Tcmp[13][14] ,
         \s_entries_Freg_Tcmp[13][13] , \s_entries_Freg_Tcmp[13][12] ,
         \s_entries_Freg_Tcmp[13][11] , \s_entries_Freg_Tcmp[13][10] ,
         \s_entries_Freg_Tcmp[13][9] , \s_entries_Freg_Tcmp[13][8] ,
         \s_entries_Freg_Tcmp[13][7] , \s_entries_Freg_Tcmp[13][6] ,
         \s_entries_Freg_Tcmp[13][5] , \s_entries_Freg_Tcmp[13][4] ,
         \s_entries_Freg_Tcmp[13][3] , \s_entries_Freg_Tcmp[13][2] ,
         \s_entries_Freg_Tcmp[13][1] , \s_entries_Freg_Tcmp[13][0] ,
         \s_entries_Freg_Tcmp[14][31] , \s_entries_Freg_Tcmp[14][30] ,
         \s_entries_Freg_Tcmp[14][29] , \s_entries_Freg_Tcmp[14][28] ,
         \s_entries_Freg_Tcmp[14][27] , \s_entries_Freg_Tcmp[14][26] ,
         \s_entries_Freg_Tcmp[14][25] , \s_entries_Freg_Tcmp[14][24] ,
         \s_entries_Freg_Tcmp[14][23] , \s_entries_Freg_Tcmp[14][22] ,
         \s_entries_Freg_Tcmp[14][21] , \s_entries_Freg_Tcmp[14][20] ,
         \s_entries_Freg_Tcmp[14][19] , \s_entries_Freg_Tcmp[14][18] ,
         \s_entries_Freg_Tcmp[14][17] , \s_entries_Freg_Tcmp[14][16] ,
         \s_entries_Freg_Tcmp[14][15] , \s_entries_Freg_Tcmp[14][14] ,
         \s_entries_Freg_Tcmp[14][13] , \s_entries_Freg_Tcmp[14][12] ,
         \s_entries_Freg_Tcmp[14][11] , \s_entries_Freg_Tcmp[14][10] ,
         \s_entries_Freg_Tcmp[14][9] , \s_entries_Freg_Tcmp[14][8] ,
         \s_entries_Freg_Tcmp[14][7] , \s_entries_Freg_Tcmp[14][6] ,
         \s_entries_Freg_Tcmp[14][5] , \s_entries_Freg_Tcmp[14][4] ,
         \s_entries_Freg_Tcmp[14][3] , \s_entries_Freg_Tcmp[14][2] ,
         \s_entries_Freg_Tcmp[14][1] , \s_entries_Freg_Tcmp[14][0] ,
         \s_entries_Freg_Tcmp[15][31] , \s_entries_Freg_Tcmp[15][30] ,
         \s_entries_Freg_Tcmp[15][29] , \s_entries_Freg_Tcmp[15][28] ,
         \s_entries_Freg_Tcmp[15][27] , \s_entries_Freg_Tcmp[15][26] ,
         \s_entries_Freg_Tcmp[15][25] , \s_entries_Freg_Tcmp[15][24] ,
         \s_entries_Freg_Tcmp[15][23] , \s_entries_Freg_Tcmp[15][22] ,
         \s_entries_Freg_Tcmp[15][21] , \s_entries_Freg_Tcmp[15][20] ,
         \s_entries_Freg_Tcmp[15][19] , \s_entries_Freg_Tcmp[15][18] ,
         \s_entries_Freg_Tcmp[15][17] , \s_entries_Freg_Tcmp[15][16] ,
         \s_entries_Freg_Tcmp[15][15] , \s_entries_Freg_Tcmp[15][14] ,
         \s_entries_Freg_Tcmp[15][13] , \s_entries_Freg_Tcmp[15][12] ,
         \s_entries_Freg_Tcmp[15][11] , \s_entries_Freg_Tcmp[15][10] ,
         \s_entries_Freg_Tcmp[15][9] , \s_entries_Freg_Tcmp[15][8] ,
         \s_entries_Freg_Tcmp[15][7] , \s_entries_Freg_Tcmp[15][6] ,
         \s_entries_Freg_Tcmp[15][5] , \s_entries_Freg_Tcmp[15][4] ,
         \s_entries_Freg_Tcmp[15][3] , \s_entries_Freg_Tcmp[15][2] ,
         \s_entries_Freg_Tcmp[15][1] , \s_entries_Freg_Tcmp[15][0] ,
         \s_entries_Freg_Tcmp[16][31] , \s_entries_Freg_Tcmp[16][30] ,
         \s_entries_Freg_Tcmp[16][29] , \s_entries_Freg_Tcmp[16][28] ,
         \s_entries_Freg_Tcmp[16][27] , \s_entries_Freg_Tcmp[16][26] ,
         \s_entries_Freg_Tcmp[16][25] , \s_entries_Freg_Tcmp[16][24] ,
         \s_entries_Freg_Tcmp[16][23] , \s_entries_Freg_Tcmp[16][22] ,
         \s_entries_Freg_Tcmp[16][21] , \s_entries_Freg_Tcmp[16][20] ,
         \s_entries_Freg_Tcmp[16][19] , \s_entries_Freg_Tcmp[16][18] ,
         \s_entries_Freg_Tcmp[16][17] , \s_entries_Freg_Tcmp[16][16] ,
         \s_entries_Freg_Tcmp[16][15] , \s_entries_Freg_Tcmp[16][14] ,
         \s_entries_Freg_Tcmp[16][13] , \s_entries_Freg_Tcmp[16][12] ,
         \s_entries_Freg_Tcmp[16][11] , \s_entries_Freg_Tcmp[16][10] ,
         \s_entries_Freg_Tcmp[16][9] , \s_entries_Freg_Tcmp[16][8] ,
         \s_entries_Freg_Tcmp[16][7] , \s_entries_Freg_Tcmp[16][6] ,
         \s_entries_Freg_Tcmp[16][5] , \s_entries_Freg_Tcmp[16][4] ,
         \s_entries_Freg_Tcmp[16][3] , \s_entries_Freg_Tcmp[16][2] ,
         \s_entries_Freg_Tcmp[16][1] , \s_entries_Freg_Tcmp[16][0] ,
         \s_entries_Freg_Tcmp[17][31] , \s_entries_Freg_Tcmp[17][30] ,
         \s_entries_Freg_Tcmp[17][29] , \s_entries_Freg_Tcmp[17][28] ,
         \s_entries_Freg_Tcmp[17][27] , \s_entries_Freg_Tcmp[17][26] ,
         \s_entries_Freg_Tcmp[17][25] , \s_entries_Freg_Tcmp[17][24] ,
         \s_entries_Freg_Tcmp[17][23] , \s_entries_Freg_Tcmp[17][22] ,
         \s_entries_Freg_Tcmp[17][21] , \s_entries_Freg_Tcmp[17][20] ,
         \s_entries_Freg_Tcmp[17][19] , \s_entries_Freg_Tcmp[17][18] ,
         \s_entries_Freg_Tcmp[17][17] , \s_entries_Freg_Tcmp[17][16] ,
         \s_entries_Freg_Tcmp[17][15] , \s_entries_Freg_Tcmp[17][14] ,
         \s_entries_Freg_Tcmp[17][13] , \s_entries_Freg_Tcmp[17][12] ,
         \s_entries_Freg_Tcmp[17][11] , \s_entries_Freg_Tcmp[17][10] ,
         \s_entries_Freg_Tcmp[17][9] , \s_entries_Freg_Tcmp[17][8] ,
         \s_entries_Freg_Tcmp[17][7] , \s_entries_Freg_Tcmp[17][6] ,
         \s_entries_Freg_Tcmp[17][5] , \s_entries_Freg_Tcmp[17][4] ,
         \s_entries_Freg_Tcmp[17][3] , \s_entries_Freg_Tcmp[17][2] ,
         \s_entries_Freg_Tcmp[17][1] , \s_entries_Freg_Tcmp[17][0] ,
         \s_entries_Freg_Tcmp[18][31] , \s_entries_Freg_Tcmp[18][30] ,
         \s_entries_Freg_Tcmp[18][29] , \s_entries_Freg_Tcmp[18][28] ,
         \s_entries_Freg_Tcmp[18][27] , \s_entries_Freg_Tcmp[18][26] ,
         \s_entries_Freg_Tcmp[18][25] , \s_entries_Freg_Tcmp[18][24] ,
         \s_entries_Freg_Tcmp[18][23] , \s_entries_Freg_Tcmp[18][22] ,
         \s_entries_Freg_Tcmp[18][21] , \s_entries_Freg_Tcmp[18][20] ,
         \s_entries_Freg_Tcmp[18][19] , \s_entries_Freg_Tcmp[18][18] ,
         \s_entries_Freg_Tcmp[18][17] , \s_entries_Freg_Tcmp[18][16] ,
         \s_entries_Freg_Tcmp[18][15] , \s_entries_Freg_Tcmp[18][14] ,
         \s_entries_Freg_Tcmp[18][13] , \s_entries_Freg_Tcmp[18][12] ,
         \s_entries_Freg_Tcmp[18][11] , \s_entries_Freg_Tcmp[18][10] ,
         \s_entries_Freg_Tcmp[18][9] , \s_entries_Freg_Tcmp[18][8] ,
         \s_entries_Freg_Tcmp[18][7] , \s_entries_Freg_Tcmp[18][6] ,
         \s_entries_Freg_Tcmp[18][5] , \s_entries_Freg_Tcmp[18][4] ,
         \s_entries_Freg_Tcmp[18][3] , \s_entries_Freg_Tcmp[18][2] ,
         \s_entries_Freg_Tcmp[18][1] , \s_entries_Freg_Tcmp[18][0] ,
         \s_entries_Freg_Tcmp[19][31] , \s_entries_Freg_Tcmp[19][30] ,
         \s_entries_Freg_Tcmp[19][29] , \s_entries_Freg_Tcmp[19][28] ,
         \s_entries_Freg_Tcmp[19][27] , \s_entries_Freg_Tcmp[19][26] ,
         \s_entries_Freg_Tcmp[19][25] , \s_entries_Freg_Tcmp[19][24] ,
         \s_entries_Freg_Tcmp[19][23] , \s_entries_Freg_Tcmp[19][22] ,
         \s_entries_Freg_Tcmp[19][21] , \s_entries_Freg_Tcmp[19][20] ,
         \s_entries_Freg_Tcmp[19][19] , \s_entries_Freg_Tcmp[19][18] ,
         \s_entries_Freg_Tcmp[19][17] , \s_entries_Freg_Tcmp[19][16] ,
         \s_entries_Freg_Tcmp[19][15] , \s_entries_Freg_Tcmp[19][14] ,
         \s_entries_Freg_Tcmp[19][13] , \s_entries_Freg_Tcmp[19][12] ,
         \s_entries_Freg_Tcmp[19][11] , \s_entries_Freg_Tcmp[19][10] ,
         \s_entries_Freg_Tcmp[19][9] , \s_entries_Freg_Tcmp[19][8] ,
         \s_entries_Freg_Tcmp[19][7] , \s_entries_Freg_Tcmp[19][6] ,
         \s_entries_Freg_Tcmp[19][5] , \s_entries_Freg_Tcmp[19][4] ,
         \s_entries_Freg_Tcmp[19][3] , \s_entries_Freg_Tcmp[19][2] ,
         \s_entries_Freg_Tcmp[19][1] , \s_entries_Freg_Tcmp[19][0] ,
         \s_entries_Freg_Tcmp[20][31] , \s_entries_Freg_Tcmp[20][30] ,
         \s_entries_Freg_Tcmp[20][29] , \s_entries_Freg_Tcmp[20][28] ,
         \s_entries_Freg_Tcmp[20][27] , \s_entries_Freg_Tcmp[20][26] ,
         \s_entries_Freg_Tcmp[20][25] , \s_entries_Freg_Tcmp[20][24] ,
         \s_entries_Freg_Tcmp[20][23] , \s_entries_Freg_Tcmp[20][22] ,
         \s_entries_Freg_Tcmp[20][21] , \s_entries_Freg_Tcmp[20][20] ,
         \s_entries_Freg_Tcmp[20][19] , \s_entries_Freg_Tcmp[20][18] ,
         \s_entries_Freg_Tcmp[20][17] , \s_entries_Freg_Tcmp[20][16] ,
         \s_entries_Freg_Tcmp[20][15] , \s_entries_Freg_Tcmp[20][14] ,
         \s_entries_Freg_Tcmp[20][13] , \s_entries_Freg_Tcmp[20][12] ,
         \s_entries_Freg_Tcmp[20][11] , \s_entries_Freg_Tcmp[20][10] ,
         \s_entries_Freg_Tcmp[20][9] , \s_entries_Freg_Tcmp[20][8] ,
         \s_entries_Freg_Tcmp[20][7] , \s_entries_Freg_Tcmp[20][6] ,
         \s_entries_Freg_Tcmp[20][5] , \s_entries_Freg_Tcmp[20][4] ,
         \s_entries_Freg_Tcmp[20][3] , \s_entries_Freg_Tcmp[20][2] ,
         \s_entries_Freg_Tcmp[20][1] , \s_entries_Freg_Tcmp[20][0] ,
         \s_entries_Freg_Tcmp[21][31] , \s_entries_Freg_Tcmp[21][30] ,
         \s_entries_Freg_Tcmp[21][29] , \s_entries_Freg_Tcmp[21][28] ,
         \s_entries_Freg_Tcmp[21][27] , \s_entries_Freg_Tcmp[21][26] ,
         \s_entries_Freg_Tcmp[21][25] , \s_entries_Freg_Tcmp[21][24] ,
         \s_entries_Freg_Tcmp[21][23] , \s_entries_Freg_Tcmp[21][22] ,
         \s_entries_Freg_Tcmp[21][21] , \s_entries_Freg_Tcmp[21][20] ,
         \s_entries_Freg_Tcmp[21][19] , \s_entries_Freg_Tcmp[21][18] ,
         \s_entries_Freg_Tcmp[21][17] , \s_entries_Freg_Tcmp[21][16] ,
         \s_entries_Freg_Tcmp[21][15] , \s_entries_Freg_Tcmp[21][14] ,
         \s_entries_Freg_Tcmp[21][13] , \s_entries_Freg_Tcmp[21][12] ,
         \s_entries_Freg_Tcmp[21][11] , \s_entries_Freg_Tcmp[21][10] ,
         \s_entries_Freg_Tcmp[21][9] , \s_entries_Freg_Tcmp[21][8] ,
         \s_entries_Freg_Tcmp[21][7] , \s_entries_Freg_Tcmp[21][6] ,
         \s_entries_Freg_Tcmp[21][5] , \s_entries_Freg_Tcmp[21][4] ,
         \s_entries_Freg_Tcmp[21][3] , \s_entries_Freg_Tcmp[21][2] ,
         \s_entries_Freg_Tcmp[21][1] , \s_entries_Freg_Tcmp[21][0] ,
         \s_entries_Freg_Tcmp[22][31] , \s_entries_Freg_Tcmp[22][30] ,
         \s_entries_Freg_Tcmp[22][29] , \s_entries_Freg_Tcmp[22][28] ,
         \s_entries_Freg_Tcmp[22][27] , \s_entries_Freg_Tcmp[22][26] ,
         \s_entries_Freg_Tcmp[22][25] , \s_entries_Freg_Tcmp[22][24] ,
         \s_entries_Freg_Tcmp[22][23] , \s_entries_Freg_Tcmp[22][22] ,
         \s_entries_Freg_Tcmp[22][21] , \s_entries_Freg_Tcmp[22][20] ,
         \s_entries_Freg_Tcmp[22][19] , \s_entries_Freg_Tcmp[22][18] ,
         \s_entries_Freg_Tcmp[22][17] , \s_entries_Freg_Tcmp[22][16] ,
         \s_entries_Freg_Tcmp[22][15] , \s_entries_Freg_Tcmp[22][14] ,
         \s_entries_Freg_Tcmp[22][13] , \s_entries_Freg_Tcmp[22][12] ,
         \s_entries_Freg_Tcmp[22][11] , \s_entries_Freg_Tcmp[22][10] ,
         \s_entries_Freg_Tcmp[22][9] , \s_entries_Freg_Tcmp[22][8] ,
         \s_entries_Freg_Tcmp[22][7] , \s_entries_Freg_Tcmp[22][6] ,
         \s_entries_Freg_Tcmp[22][5] , \s_entries_Freg_Tcmp[22][4] ,
         \s_entries_Freg_Tcmp[22][3] , \s_entries_Freg_Tcmp[22][2] ,
         \s_entries_Freg_Tcmp[22][1] , \s_entries_Freg_Tcmp[22][0] ,
         \s_entries_Freg_Tcmp[23][31] , \s_entries_Freg_Tcmp[23][30] ,
         \s_entries_Freg_Tcmp[23][29] , \s_entries_Freg_Tcmp[23][28] ,
         \s_entries_Freg_Tcmp[23][27] , \s_entries_Freg_Tcmp[23][26] ,
         \s_entries_Freg_Tcmp[23][25] , \s_entries_Freg_Tcmp[23][24] ,
         \s_entries_Freg_Tcmp[23][23] , \s_entries_Freg_Tcmp[23][22] ,
         \s_entries_Freg_Tcmp[23][21] , \s_entries_Freg_Tcmp[23][20] ,
         \s_entries_Freg_Tcmp[23][19] , \s_entries_Freg_Tcmp[23][18] ,
         \s_entries_Freg_Tcmp[23][17] , \s_entries_Freg_Tcmp[23][16] ,
         \s_entries_Freg_Tcmp[23][15] , \s_entries_Freg_Tcmp[23][14] ,
         \s_entries_Freg_Tcmp[23][13] , \s_entries_Freg_Tcmp[23][12] ,
         \s_entries_Freg_Tcmp[23][11] , \s_entries_Freg_Tcmp[23][10] ,
         \s_entries_Freg_Tcmp[23][9] , \s_entries_Freg_Tcmp[23][8] ,
         \s_entries_Freg_Tcmp[23][7] , \s_entries_Freg_Tcmp[23][6] ,
         \s_entries_Freg_Tcmp[23][5] , \s_entries_Freg_Tcmp[23][4] ,
         \s_entries_Freg_Tcmp[23][3] , \s_entries_Freg_Tcmp[23][2] ,
         \s_entries_Freg_Tcmp[23][1] , \s_entries_Freg_Tcmp[23][0] ,
         \s_entries_Freg_Tcmp[24][31] , \s_entries_Freg_Tcmp[24][30] ,
         \s_entries_Freg_Tcmp[24][29] , \s_entries_Freg_Tcmp[24][28] ,
         \s_entries_Freg_Tcmp[24][27] , \s_entries_Freg_Tcmp[24][26] ,
         \s_entries_Freg_Tcmp[24][25] , \s_entries_Freg_Tcmp[24][24] ,
         \s_entries_Freg_Tcmp[24][23] , \s_entries_Freg_Tcmp[24][22] ,
         \s_entries_Freg_Tcmp[24][21] , \s_entries_Freg_Tcmp[24][20] ,
         \s_entries_Freg_Tcmp[24][19] , \s_entries_Freg_Tcmp[24][18] ,
         \s_entries_Freg_Tcmp[24][17] , \s_entries_Freg_Tcmp[24][16] ,
         \s_entries_Freg_Tcmp[24][15] , \s_entries_Freg_Tcmp[24][14] ,
         \s_entries_Freg_Tcmp[24][13] , \s_entries_Freg_Tcmp[24][12] ,
         \s_entries_Freg_Tcmp[24][11] , \s_entries_Freg_Tcmp[24][10] ,
         \s_entries_Freg_Tcmp[24][9] , \s_entries_Freg_Tcmp[24][8] ,
         \s_entries_Freg_Tcmp[24][7] , \s_entries_Freg_Tcmp[24][6] ,
         \s_entries_Freg_Tcmp[24][5] , \s_entries_Freg_Tcmp[24][4] ,
         \s_entries_Freg_Tcmp[24][3] , \s_entries_Freg_Tcmp[24][2] ,
         \s_entries_Freg_Tcmp[24][1] , \s_entries_Freg_Tcmp[24][0] ,
         \s_entries_Freg_Tcmp[25][31] , \s_entries_Freg_Tcmp[25][30] ,
         \s_entries_Freg_Tcmp[25][29] , \s_entries_Freg_Tcmp[25][28] ,
         \s_entries_Freg_Tcmp[25][27] , \s_entries_Freg_Tcmp[25][26] ,
         \s_entries_Freg_Tcmp[25][25] , \s_entries_Freg_Tcmp[25][24] ,
         \s_entries_Freg_Tcmp[25][23] , \s_entries_Freg_Tcmp[25][22] ,
         \s_entries_Freg_Tcmp[25][21] , \s_entries_Freg_Tcmp[25][20] ,
         \s_entries_Freg_Tcmp[25][19] , \s_entries_Freg_Tcmp[25][18] ,
         \s_entries_Freg_Tcmp[25][17] , \s_entries_Freg_Tcmp[25][16] ,
         \s_entries_Freg_Tcmp[25][15] , \s_entries_Freg_Tcmp[25][14] ,
         \s_entries_Freg_Tcmp[25][13] , \s_entries_Freg_Tcmp[25][12] ,
         \s_entries_Freg_Tcmp[25][11] , \s_entries_Freg_Tcmp[25][10] ,
         \s_entries_Freg_Tcmp[25][9] , \s_entries_Freg_Tcmp[25][8] ,
         \s_entries_Freg_Tcmp[25][7] , \s_entries_Freg_Tcmp[25][6] ,
         \s_entries_Freg_Tcmp[25][5] , \s_entries_Freg_Tcmp[25][4] ,
         \s_entries_Freg_Tcmp[25][3] , \s_entries_Freg_Tcmp[25][2] ,
         \s_entries_Freg_Tcmp[25][1] , \s_entries_Freg_Tcmp[25][0] ,
         \s_entries_Freg_Tcmp[26][31] , \s_entries_Freg_Tcmp[26][30] ,
         \s_entries_Freg_Tcmp[26][29] , \s_entries_Freg_Tcmp[26][28] ,
         \s_entries_Freg_Tcmp[26][27] , \s_entries_Freg_Tcmp[26][26] ,
         \s_entries_Freg_Tcmp[26][25] , \s_entries_Freg_Tcmp[26][24] ,
         \s_entries_Freg_Tcmp[26][23] , \s_entries_Freg_Tcmp[26][22] ,
         \s_entries_Freg_Tcmp[26][21] , \s_entries_Freg_Tcmp[26][20] ,
         \s_entries_Freg_Tcmp[26][19] , \s_entries_Freg_Tcmp[26][18] ,
         \s_entries_Freg_Tcmp[26][17] , \s_entries_Freg_Tcmp[26][16] ,
         \s_entries_Freg_Tcmp[26][15] , \s_entries_Freg_Tcmp[26][14] ,
         \s_entries_Freg_Tcmp[26][13] , \s_entries_Freg_Tcmp[26][12] ,
         \s_entries_Freg_Tcmp[26][11] , \s_entries_Freg_Tcmp[26][10] ,
         \s_entries_Freg_Tcmp[26][9] , \s_entries_Freg_Tcmp[26][8] ,
         \s_entries_Freg_Tcmp[26][7] , \s_entries_Freg_Tcmp[26][6] ,
         \s_entries_Freg_Tcmp[26][5] , \s_entries_Freg_Tcmp[26][4] ,
         \s_entries_Freg_Tcmp[26][3] , \s_entries_Freg_Tcmp[26][2] ,
         \s_entries_Freg_Tcmp[26][1] , \s_entries_Freg_Tcmp[26][0] ,
         \s_entries_Freg_Tcmp[27][31] , \s_entries_Freg_Tcmp[27][30] ,
         \s_entries_Freg_Tcmp[27][29] , \s_entries_Freg_Tcmp[27][28] ,
         \s_entries_Freg_Tcmp[27][27] , \s_entries_Freg_Tcmp[27][26] ,
         \s_entries_Freg_Tcmp[27][25] , \s_entries_Freg_Tcmp[27][24] ,
         \s_entries_Freg_Tcmp[27][23] , \s_entries_Freg_Tcmp[27][22] ,
         \s_entries_Freg_Tcmp[27][21] , \s_entries_Freg_Tcmp[27][20] ,
         \s_entries_Freg_Tcmp[27][19] , \s_entries_Freg_Tcmp[27][18] ,
         \s_entries_Freg_Tcmp[27][17] , \s_entries_Freg_Tcmp[27][16] ,
         \s_entries_Freg_Tcmp[27][15] , \s_entries_Freg_Tcmp[27][14] ,
         \s_entries_Freg_Tcmp[27][13] , \s_entries_Freg_Tcmp[27][12] ,
         \s_entries_Freg_Tcmp[27][11] , \s_entries_Freg_Tcmp[27][10] ,
         \s_entries_Freg_Tcmp[27][9] , \s_entries_Freg_Tcmp[27][8] ,
         \s_entries_Freg_Tcmp[27][7] , \s_entries_Freg_Tcmp[27][6] ,
         \s_entries_Freg_Tcmp[27][5] , \s_entries_Freg_Tcmp[27][4] ,
         \s_entries_Freg_Tcmp[27][3] , \s_entries_Freg_Tcmp[27][2] ,
         \s_entries_Freg_Tcmp[27][1] , \s_entries_Freg_Tcmp[27][0] ,
         \s_entries_Freg_Tcmp[28][31] , \s_entries_Freg_Tcmp[28][30] ,
         \s_entries_Freg_Tcmp[28][29] , \s_entries_Freg_Tcmp[28][28] ,
         \s_entries_Freg_Tcmp[28][27] , \s_entries_Freg_Tcmp[28][26] ,
         \s_entries_Freg_Tcmp[28][25] , \s_entries_Freg_Tcmp[28][24] ,
         \s_entries_Freg_Tcmp[28][23] , \s_entries_Freg_Tcmp[28][22] ,
         \s_entries_Freg_Tcmp[28][21] , \s_entries_Freg_Tcmp[28][20] ,
         \s_entries_Freg_Tcmp[28][19] , \s_entries_Freg_Tcmp[28][18] ,
         \s_entries_Freg_Tcmp[28][17] , \s_entries_Freg_Tcmp[28][16] ,
         \s_entries_Freg_Tcmp[28][15] , \s_entries_Freg_Tcmp[28][14] ,
         \s_entries_Freg_Tcmp[28][13] , \s_entries_Freg_Tcmp[28][12] ,
         \s_entries_Freg_Tcmp[28][11] , \s_entries_Freg_Tcmp[28][10] ,
         \s_entries_Freg_Tcmp[28][9] , \s_entries_Freg_Tcmp[28][8] ,
         \s_entries_Freg_Tcmp[28][7] , \s_entries_Freg_Tcmp[28][6] ,
         \s_entries_Freg_Tcmp[28][5] , \s_entries_Freg_Tcmp[28][4] ,
         \s_entries_Freg_Tcmp[28][3] , \s_entries_Freg_Tcmp[28][2] ,
         \s_entries_Freg_Tcmp[28][1] , \s_entries_Freg_Tcmp[28][0] ,
         \s_entries_Freg_Tcmp[29][31] , \s_entries_Freg_Tcmp[29][30] ,
         \s_entries_Freg_Tcmp[29][29] , \s_entries_Freg_Tcmp[29][28] ,
         \s_entries_Freg_Tcmp[29][27] , \s_entries_Freg_Tcmp[29][26] ,
         \s_entries_Freg_Tcmp[29][25] , \s_entries_Freg_Tcmp[29][24] ,
         \s_entries_Freg_Tcmp[29][23] , \s_entries_Freg_Tcmp[29][22] ,
         \s_entries_Freg_Tcmp[29][21] , \s_entries_Freg_Tcmp[29][20] ,
         \s_entries_Freg_Tcmp[29][19] , \s_entries_Freg_Tcmp[29][18] ,
         \s_entries_Freg_Tcmp[29][17] , \s_entries_Freg_Tcmp[29][16] ,
         \s_entries_Freg_Tcmp[29][15] , \s_entries_Freg_Tcmp[29][14] ,
         \s_entries_Freg_Tcmp[29][13] , \s_entries_Freg_Tcmp[29][12] ,
         \s_entries_Freg_Tcmp[29][11] , \s_entries_Freg_Tcmp[29][10] ,
         \s_entries_Freg_Tcmp[29][9] , \s_entries_Freg_Tcmp[29][8] ,
         \s_entries_Freg_Tcmp[29][7] , \s_entries_Freg_Tcmp[29][6] ,
         \s_entries_Freg_Tcmp[29][5] , \s_entries_Freg_Tcmp[29][4] ,
         \s_entries_Freg_Tcmp[29][3] , \s_entries_Freg_Tcmp[29][2] ,
         \s_entries_Freg_Tcmp[29][1] , \s_entries_Freg_Tcmp[29][0] ,
         \s_entries_Freg_Tcmp[30][31] , \s_entries_Freg_Tcmp[30][30] ,
         \s_entries_Freg_Tcmp[30][29] , \s_entries_Freg_Tcmp[30][28] ,
         \s_entries_Freg_Tcmp[30][27] , \s_entries_Freg_Tcmp[30][26] ,
         \s_entries_Freg_Tcmp[30][25] , \s_entries_Freg_Tcmp[30][24] ,
         \s_entries_Freg_Tcmp[30][23] , \s_entries_Freg_Tcmp[30][22] ,
         \s_entries_Freg_Tcmp[30][21] , \s_entries_Freg_Tcmp[30][20] ,
         \s_entries_Freg_Tcmp[30][19] , \s_entries_Freg_Tcmp[30][18] ,
         \s_entries_Freg_Tcmp[30][17] , \s_entries_Freg_Tcmp[30][16] ,
         \s_entries_Freg_Tcmp[30][15] , \s_entries_Freg_Tcmp[30][14] ,
         \s_entries_Freg_Tcmp[30][13] , \s_entries_Freg_Tcmp[30][12] ,
         \s_entries_Freg_Tcmp[30][11] , \s_entries_Freg_Tcmp[30][10] ,
         \s_entries_Freg_Tcmp[30][9] , \s_entries_Freg_Tcmp[30][8] ,
         \s_entries_Freg_Tcmp[30][7] , \s_entries_Freg_Tcmp[30][6] ,
         \s_entries_Freg_Tcmp[30][5] , \s_entries_Freg_Tcmp[30][4] ,
         \s_entries_Freg_Tcmp[30][3] , \s_entries_Freg_Tcmp[30][2] ,
         \s_entries_Freg_Tcmp[30][1] , \s_entries_Freg_Tcmp[30][0] ,
         \s_entries_Freg_Tcmp[31][31] , \s_entries_Freg_Tcmp[31][30] ,
         \s_entries_Freg_Tcmp[31][29] , \s_entries_Freg_Tcmp[31][28] ,
         \s_entries_Freg_Tcmp[31][27] , \s_entries_Freg_Tcmp[31][26] ,
         \s_entries_Freg_Tcmp[31][25] , \s_entries_Freg_Tcmp[31][24] ,
         \s_entries_Freg_Tcmp[31][23] , \s_entries_Freg_Tcmp[31][22] ,
         \s_entries_Freg_Tcmp[31][21] , \s_entries_Freg_Tcmp[31][20] ,
         \s_entries_Freg_Tcmp[31][19] , \s_entries_Freg_Tcmp[31][18] ,
         \s_entries_Freg_Tcmp[31][17] , \s_entries_Freg_Tcmp[31][16] ,
         \s_entries_Freg_Tcmp[31][15] , \s_entries_Freg_Tcmp[31][14] ,
         \s_entries_Freg_Tcmp[31][13] , \s_entries_Freg_Tcmp[31][12] ,
         \s_entries_Freg_Tcmp[31][11] , \s_entries_Freg_Tcmp[31][10] ,
         \s_entries_Freg_Tcmp[31][9] , \s_entries_Freg_Tcmp[31][8] ,
         \s_entries_Freg_Tcmp[31][7] , \s_entries_Freg_Tcmp[31][6] ,
         \s_entries_Freg_Tcmp[31][5] , \s_entries_Freg_Tcmp[31][4] ,
         \s_entries_Freg_Tcmp[31][3] , \s_entries_Freg_Tcmp[31][2] ,
         \s_entries_Freg_Tcmp[31][1] , \s_entries_Freg_Tcmp[31][0] ,
         s_HIT_miss, \s_mux_signals[0][0][31] , \s_mux_signals[0][0][30] ,
         \s_mux_signals[0][0][29] , \s_mux_signals[0][0][28] ,
         \s_mux_signals[0][0][27] , \s_mux_signals[0][0][26] ,
         \s_mux_signals[0][0][25] , \s_mux_signals[0][0][24] ,
         \s_mux_signals[0][0][23] , \s_mux_signals[0][0][22] ,
         \s_mux_signals[0][0][21] , \s_mux_signals[0][0][20] ,
         \s_mux_signals[0][0][19] , \s_mux_signals[0][0][18] ,
         \s_mux_signals[0][0][17] , \s_mux_signals[0][0][16] ,
         \s_mux_signals[0][0][15] , \s_mux_signals[0][0][14] ,
         \s_mux_signals[0][0][13] , \s_mux_signals[0][0][12] ,
         \s_mux_signals[0][0][11] , \s_mux_signals[0][0][10] ,
         \s_mux_signals[0][0][9] , \s_mux_signals[0][0][8] ,
         \s_mux_signals[0][0][7] , \s_mux_signals[0][0][6] ,
         \s_mux_signals[0][0][5] , \s_mux_signals[0][0][4] ,
         \s_mux_signals[0][0][3] , \s_mux_signals[0][0][2] ,
         \s_mux_signals[0][0][1] , \s_mux_signals[0][0][0] ,
         \s_mux_signals[0][1][31] , \s_mux_signals[0][1][30] ,
         \s_mux_signals[0][1][29] , \s_mux_signals[0][1][28] ,
         \s_mux_signals[0][1][27] , \s_mux_signals[0][1][26] ,
         \s_mux_signals[0][1][25] , \s_mux_signals[0][1][24] ,
         \s_mux_signals[0][1][23] , \s_mux_signals[0][1][22] ,
         \s_mux_signals[0][1][21] , \s_mux_signals[0][1][20] ,
         \s_mux_signals[0][1][19] , \s_mux_signals[0][1][18] ,
         \s_mux_signals[0][1][17] , \s_mux_signals[0][1][16] ,
         \s_mux_signals[0][1][15] , \s_mux_signals[0][1][14] ,
         \s_mux_signals[0][1][13] , \s_mux_signals[0][1][12] ,
         \s_mux_signals[0][1][11] , \s_mux_signals[0][1][10] ,
         \s_mux_signals[0][1][9] , \s_mux_signals[0][1][8] ,
         \s_mux_signals[0][1][7] , \s_mux_signals[0][1][6] ,
         \s_mux_signals[0][1][5] , \s_mux_signals[0][1][4] ,
         \s_mux_signals[0][1][3] , \s_mux_signals[0][1][2] ,
         \s_mux_signals[0][1][1] , \s_mux_signals[0][1][0] ,
         \s_mux_signals[0][2][31] , \s_mux_signals[0][2][30] ,
         \s_mux_signals[0][2][29] , \s_mux_signals[0][2][28] ,
         \s_mux_signals[0][2][27] , \s_mux_signals[0][2][26] ,
         \s_mux_signals[0][2][25] , \s_mux_signals[0][2][24] ,
         \s_mux_signals[0][2][23] , \s_mux_signals[0][2][22] ,
         \s_mux_signals[0][2][21] , \s_mux_signals[0][2][20] ,
         \s_mux_signals[0][2][19] , \s_mux_signals[0][2][18] ,
         \s_mux_signals[0][2][17] , \s_mux_signals[0][2][16] ,
         \s_mux_signals[0][2][15] , \s_mux_signals[0][2][14] ,
         \s_mux_signals[0][2][13] , \s_mux_signals[0][2][12] ,
         \s_mux_signals[0][2][11] , \s_mux_signals[0][2][10] ,
         \s_mux_signals[0][2][9] , \s_mux_signals[0][2][8] ,
         \s_mux_signals[0][2][7] , \s_mux_signals[0][2][6] ,
         \s_mux_signals[0][2][5] , \s_mux_signals[0][2][4] ,
         \s_mux_signals[0][2][3] , \s_mux_signals[0][2][2] ,
         \s_mux_signals[0][2][1] , \s_mux_signals[0][2][0] ,
         \s_mux_signals[0][3][31] , \s_mux_signals[0][3][30] ,
         \s_mux_signals[0][3][29] , \s_mux_signals[0][3][28] ,
         \s_mux_signals[0][3][27] , \s_mux_signals[0][3][26] ,
         \s_mux_signals[0][3][25] , \s_mux_signals[0][3][24] ,
         \s_mux_signals[0][3][23] , \s_mux_signals[0][3][22] ,
         \s_mux_signals[0][3][21] , \s_mux_signals[0][3][20] ,
         \s_mux_signals[0][3][19] , \s_mux_signals[0][3][18] ,
         \s_mux_signals[0][3][17] , \s_mux_signals[0][3][16] ,
         \s_mux_signals[0][3][15] , \s_mux_signals[0][3][14] ,
         \s_mux_signals[0][3][13] , \s_mux_signals[0][3][12] ,
         \s_mux_signals[0][3][11] , \s_mux_signals[0][3][10] ,
         \s_mux_signals[0][3][9] , \s_mux_signals[0][3][8] ,
         \s_mux_signals[0][3][7] , \s_mux_signals[0][3][6] ,
         \s_mux_signals[0][3][5] , \s_mux_signals[0][3][4] ,
         \s_mux_signals[0][3][3] , \s_mux_signals[0][3][2] ,
         \s_mux_signals[0][3][1] , \s_mux_signals[0][3][0] ,
         \s_mux_signals[0][4][31] , \s_mux_signals[0][4][30] ,
         \s_mux_signals[0][4][29] , \s_mux_signals[0][4][28] ,
         \s_mux_signals[0][4][27] , \s_mux_signals[0][4][26] ,
         \s_mux_signals[0][4][25] , \s_mux_signals[0][4][24] ,
         \s_mux_signals[0][4][23] , \s_mux_signals[0][4][22] ,
         \s_mux_signals[0][4][21] , \s_mux_signals[0][4][20] ,
         \s_mux_signals[0][4][19] , \s_mux_signals[0][4][18] ,
         \s_mux_signals[0][4][17] , \s_mux_signals[0][4][16] ,
         \s_mux_signals[0][4][15] , \s_mux_signals[0][4][14] ,
         \s_mux_signals[0][4][13] , \s_mux_signals[0][4][12] ,
         \s_mux_signals[0][4][11] , \s_mux_signals[0][4][10] ,
         \s_mux_signals[0][4][9] , \s_mux_signals[0][4][8] ,
         \s_mux_signals[0][4][7] , \s_mux_signals[0][4][6] ,
         \s_mux_signals[0][4][5] , \s_mux_signals[0][4][4] ,
         \s_mux_signals[0][4][3] , \s_mux_signals[0][4][2] ,
         \s_mux_signals[0][4][1] , \s_mux_signals[0][4][0] ,
         \s_mux_signals[0][5][31] , \s_mux_signals[0][5][30] ,
         \s_mux_signals[0][5][29] , \s_mux_signals[0][5][28] ,
         \s_mux_signals[0][5][27] , \s_mux_signals[0][5][26] ,
         \s_mux_signals[0][5][25] , \s_mux_signals[0][5][24] ,
         \s_mux_signals[0][5][23] , \s_mux_signals[0][5][22] ,
         \s_mux_signals[0][5][21] , \s_mux_signals[0][5][20] ,
         \s_mux_signals[0][5][19] , \s_mux_signals[0][5][18] ,
         \s_mux_signals[0][5][17] , \s_mux_signals[0][5][16] ,
         \s_mux_signals[0][5][15] , \s_mux_signals[0][5][14] ,
         \s_mux_signals[0][5][13] , \s_mux_signals[0][5][12] ,
         \s_mux_signals[0][5][11] , \s_mux_signals[0][5][10] ,
         \s_mux_signals[0][5][9] , \s_mux_signals[0][5][8] ,
         \s_mux_signals[0][5][7] , \s_mux_signals[0][5][6] ,
         \s_mux_signals[0][5][5] , \s_mux_signals[0][5][4] ,
         \s_mux_signals[0][5][3] , \s_mux_signals[0][5][2] ,
         \s_mux_signals[0][5][1] , \s_mux_signals[0][5][0] ,
         \s_mux_signals[0][6][31] , \s_mux_signals[0][6][30] ,
         \s_mux_signals[0][6][29] , \s_mux_signals[0][6][28] ,
         \s_mux_signals[0][6][27] , \s_mux_signals[0][6][26] ,
         \s_mux_signals[0][6][25] , \s_mux_signals[0][6][24] ,
         \s_mux_signals[0][6][23] , \s_mux_signals[0][6][22] ,
         \s_mux_signals[0][6][21] , \s_mux_signals[0][6][20] ,
         \s_mux_signals[0][6][19] , \s_mux_signals[0][6][18] ,
         \s_mux_signals[0][6][17] , \s_mux_signals[0][6][16] ,
         \s_mux_signals[0][6][15] , \s_mux_signals[0][6][14] ,
         \s_mux_signals[0][6][13] , \s_mux_signals[0][6][12] ,
         \s_mux_signals[0][6][11] , \s_mux_signals[0][6][10] ,
         \s_mux_signals[0][6][9] , \s_mux_signals[0][6][8] ,
         \s_mux_signals[0][6][7] , \s_mux_signals[0][6][6] ,
         \s_mux_signals[0][6][5] , \s_mux_signals[0][6][4] ,
         \s_mux_signals[0][6][3] , \s_mux_signals[0][6][2] ,
         \s_mux_signals[0][6][1] , \s_mux_signals[0][6][0] ,
         \s_mux_signals[0][7][31] , \s_mux_signals[0][7][30] ,
         \s_mux_signals[0][7][29] , \s_mux_signals[0][7][28] ,
         \s_mux_signals[0][7][27] , \s_mux_signals[0][7][26] ,
         \s_mux_signals[0][7][25] , \s_mux_signals[0][7][24] ,
         \s_mux_signals[0][7][23] , \s_mux_signals[0][7][22] ,
         \s_mux_signals[0][7][21] , \s_mux_signals[0][7][20] ,
         \s_mux_signals[0][7][19] , \s_mux_signals[0][7][18] ,
         \s_mux_signals[0][7][17] , \s_mux_signals[0][7][16] ,
         \s_mux_signals[0][7][15] , \s_mux_signals[0][7][14] ,
         \s_mux_signals[0][7][13] , \s_mux_signals[0][7][12] ,
         \s_mux_signals[0][7][11] , \s_mux_signals[0][7][10] ,
         \s_mux_signals[0][7][9] , \s_mux_signals[0][7][8] ,
         \s_mux_signals[0][7][7] , \s_mux_signals[0][7][6] ,
         \s_mux_signals[0][7][5] , \s_mux_signals[0][7][4] ,
         \s_mux_signals[0][7][3] , \s_mux_signals[0][7][2] ,
         \s_mux_signals[0][7][1] , \s_mux_signals[0][7][0] ,
         \s_mux_signals[0][8][31] , \s_mux_signals[0][8][30] ,
         \s_mux_signals[0][8][29] , \s_mux_signals[0][8][28] ,
         \s_mux_signals[0][8][27] , \s_mux_signals[0][8][26] ,
         \s_mux_signals[0][8][25] , \s_mux_signals[0][8][24] ,
         \s_mux_signals[0][8][23] , \s_mux_signals[0][8][22] ,
         \s_mux_signals[0][8][21] , \s_mux_signals[0][8][20] ,
         \s_mux_signals[0][8][19] , \s_mux_signals[0][8][18] ,
         \s_mux_signals[0][8][17] , \s_mux_signals[0][8][16] ,
         \s_mux_signals[0][8][15] , \s_mux_signals[0][8][14] ,
         \s_mux_signals[0][8][13] , \s_mux_signals[0][8][12] ,
         \s_mux_signals[0][8][11] , \s_mux_signals[0][8][10] ,
         \s_mux_signals[0][8][9] , \s_mux_signals[0][8][8] ,
         \s_mux_signals[0][8][7] , \s_mux_signals[0][8][6] ,
         \s_mux_signals[0][8][5] , \s_mux_signals[0][8][4] ,
         \s_mux_signals[0][8][3] , \s_mux_signals[0][8][2] ,
         \s_mux_signals[0][8][1] , \s_mux_signals[0][8][0] ,
         \s_mux_signals[0][9][31] , \s_mux_signals[0][9][30] ,
         \s_mux_signals[0][9][29] , \s_mux_signals[0][9][28] ,
         \s_mux_signals[0][9][27] , \s_mux_signals[0][9][26] ,
         \s_mux_signals[0][9][25] , \s_mux_signals[0][9][24] ,
         \s_mux_signals[0][9][23] , \s_mux_signals[0][9][22] ,
         \s_mux_signals[0][9][21] , \s_mux_signals[0][9][20] ,
         \s_mux_signals[0][9][19] , \s_mux_signals[0][9][18] ,
         \s_mux_signals[0][9][17] , \s_mux_signals[0][9][16] ,
         \s_mux_signals[0][9][15] , \s_mux_signals[0][9][14] ,
         \s_mux_signals[0][9][13] , \s_mux_signals[0][9][12] ,
         \s_mux_signals[0][9][11] , \s_mux_signals[0][9][10] ,
         \s_mux_signals[0][9][9] , \s_mux_signals[0][9][8] ,
         \s_mux_signals[0][9][7] , \s_mux_signals[0][9][6] ,
         \s_mux_signals[0][9][5] , \s_mux_signals[0][9][4] ,
         \s_mux_signals[0][9][3] , \s_mux_signals[0][9][2] ,
         \s_mux_signals[0][9][1] , \s_mux_signals[0][9][0] ,
         \s_mux_signals[0][10][31] , \s_mux_signals[0][10][30] ,
         \s_mux_signals[0][10][29] , \s_mux_signals[0][10][28] ,
         \s_mux_signals[0][10][27] , \s_mux_signals[0][10][26] ,
         \s_mux_signals[0][10][25] , \s_mux_signals[0][10][24] ,
         \s_mux_signals[0][10][23] , \s_mux_signals[0][10][22] ,
         \s_mux_signals[0][10][21] , \s_mux_signals[0][10][20] ,
         \s_mux_signals[0][10][19] , \s_mux_signals[0][10][18] ,
         \s_mux_signals[0][10][17] , \s_mux_signals[0][10][16] ,
         \s_mux_signals[0][10][15] , \s_mux_signals[0][10][14] ,
         \s_mux_signals[0][10][13] , \s_mux_signals[0][10][12] ,
         \s_mux_signals[0][10][11] , \s_mux_signals[0][10][10] ,
         \s_mux_signals[0][10][9] , \s_mux_signals[0][10][8] ,
         \s_mux_signals[0][10][7] , \s_mux_signals[0][10][6] ,
         \s_mux_signals[0][10][5] , \s_mux_signals[0][10][4] ,
         \s_mux_signals[0][10][3] , \s_mux_signals[0][10][2] ,
         \s_mux_signals[0][10][1] , \s_mux_signals[0][10][0] ,
         \s_mux_signals[0][11][31] , \s_mux_signals[0][11][30] ,
         \s_mux_signals[0][11][29] , \s_mux_signals[0][11][28] ,
         \s_mux_signals[0][11][27] , \s_mux_signals[0][11][26] ,
         \s_mux_signals[0][11][25] , \s_mux_signals[0][11][24] ,
         \s_mux_signals[0][11][23] , \s_mux_signals[0][11][22] ,
         \s_mux_signals[0][11][21] , \s_mux_signals[0][11][20] ,
         \s_mux_signals[0][11][19] , \s_mux_signals[0][11][18] ,
         \s_mux_signals[0][11][17] , \s_mux_signals[0][11][16] ,
         \s_mux_signals[0][11][15] , \s_mux_signals[0][11][14] ,
         \s_mux_signals[0][11][13] , \s_mux_signals[0][11][12] ,
         \s_mux_signals[0][11][11] , \s_mux_signals[0][11][10] ,
         \s_mux_signals[0][11][9] , \s_mux_signals[0][11][8] ,
         \s_mux_signals[0][11][7] , \s_mux_signals[0][11][6] ,
         \s_mux_signals[0][11][5] , \s_mux_signals[0][11][4] ,
         \s_mux_signals[0][11][3] , \s_mux_signals[0][11][2] ,
         \s_mux_signals[0][11][1] , \s_mux_signals[0][11][0] ,
         \s_mux_signals[0][12][31] , \s_mux_signals[0][12][30] ,
         \s_mux_signals[0][12][29] , \s_mux_signals[0][12][28] ,
         \s_mux_signals[0][12][27] , \s_mux_signals[0][12][26] ,
         \s_mux_signals[0][12][25] , \s_mux_signals[0][12][24] ,
         \s_mux_signals[0][12][23] , \s_mux_signals[0][12][22] ,
         \s_mux_signals[0][12][21] , \s_mux_signals[0][12][20] ,
         \s_mux_signals[0][12][19] , \s_mux_signals[0][12][18] ,
         \s_mux_signals[0][12][17] , \s_mux_signals[0][12][16] ,
         \s_mux_signals[0][12][15] , \s_mux_signals[0][12][14] ,
         \s_mux_signals[0][12][13] , \s_mux_signals[0][12][12] ,
         \s_mux_signals[0][12][11] , \s_mux_signals[0][12][10] ,
         \s_mux_signals[0][12][9] , \s_mux_signals[0][12][8] ,
         \s_mux_signals[0][12][7] , \s_mux_signals[0][12][6] ,
         \s_mux_signals[0][12][5] , \s_mux_signals[0][12][4] ,
         \s_mux_signals[0][12][3] , \s_mux_signals[0][12][2] ,
         \s_mux_signals[0][12][1] , \s_mux_signals[0][12][0] ,
         \s_mux_signals[0][13][31] , \s_mux_signals[0][13][30] ,
         \s_mux_signals[0][13][29] , \s_mux_signals[0][13][28] ,
         \s_mux_signals[0][13][27] , \s_mux_signals[0][13][26] ,
         \s_mux_signals[0][13][25] , \s_mux_signals[0][13][24] ,
         \s_mux_signals[0][13][23] , \s_mux_signals[0][13][22] ,
         \s_mux_signals[0][13][21] , \s_mux_signals[0][13][20] ,
         \s_mux_signals[0][13][19] , \s_mux_signals[0][13][18] ,
         \s_mux_signals[0][13][17] , \s_mux_signals[0][13][16] ,
         \s_mux_signals[0][13][15] , \s_mux_signals[0][13][14] ,
         \s_mux_signals[0][13][13] , \s_mux_signals[0][13][12] ,
         \s_mux_signals[0][13][11] , \s_mux_signals[0][13][10] ,
         \s_mux_signals[0][13][9] , \s_mux_signals[0][13][8] ,
         \s_mux_signals[0][13][7] , \s_mux_signals[0][13][6] ,
         \s_mux_signals[0][13][5] , \s_mux_signals[0][13][4] ,
         \s_mux_signals[0][13][3] , \s_mux_signals[0][13][2] ,
         \s_mux_signals[0][13][1] , \s_mux_signals[0][13][0] ,
         \s_mux_signals[0][14][31] , \s_mux_signals[0][14][30] ,
         \s_mux_signals[0][14][29] , \s_mux_signals[0][14][28] ,
         \s_mux_signals[0][14][27] , \s_mux_signals[0][14][26] ,
         \s_mux_signals[0][14][25] , \s_mux_signals[0][14][24] ,
         \s_mux_signals[0][14][23] , \s_mux_signals[0][14][22] ,
         \s_mux_signals[0][14][21] , \s_mux_signals[0][14][20] ,
         \s_mux_signals[0][14][19] , \s_mux_signals[0][14][18] ,
         \s_mux_signals[0][14][17] , \s_mux_signals[0][14][16] ,
         \s_mux_signals[0][14][15] , \s_mux_signals[0][14][14] ,
         \s_mux_signals[0][14][13] , \s_mux_signals[0][14][12] ,
         \s_mux_signals[0][14][11] , \s_mux_signals[0][14][10] ,
         \s_mux_signals[0][14][9] , \s_mux_signals[0][14][8] ,
         \s_mux_signals[0][14][7] , \s_mux_signals[0][14][6] ,
         \s_mux_signals[0][14][5] , \s_mux_signals[0][14][4] ,
         \s_mux_signals[0][14][3] , \s_mux_signals[0][14][2] ,
         \s_mux_signals[0][14][1] , \s_mux_signals[0][14][0] ,
         \s_mux_signals[0][15][31] , \s_mux_signals[0][15][30] ,
         \s_mux_signals[0][15][29] , \s_mux_signals[0][15][28] ,
         \s_mux_signals[0][15][27] , \s_mux_signals[0][15][26] ,
         \s_mux_signals[0][15][25] , \s_mux_signals[0][15][24] ,
         \s_mux_signals[0][15][23] , \s_mux_signals[0][15][22] ,
         \s_mux_signals[0][15][21] , \s_mux_signals[0][15][20] ,
         \s_mux_signals[0][15][19] , \s_mux_signals[0][15][18] ,
         \s_mux_signals[0][15][17] , \s_mux_signals[0][15][16] ,
         \s_mux_signals[0][15][15] , \s_mux_signals[0][15][14] ,
         \s_mux_signals[0][15][13] , \s_mux_signals[0][15][12] ,
         \s_mux_signals[0][15][11] , \s_mux_signals[0][15][10] ,
         \s_mux_signals[0][15][9] , \s_mux_signals[0][15][8] ,
         \s_mux_signals[0][15][7] , \s_mux_signals[0][15][6] ,
         \s_mux_signals[0][15][5] , \s_mux_signals[0][15][4] ,
         \s_mux_signals[0][15][3] , \s_mux_signals[0][15][2] ,
         \s_mux_signals[0][15][1] , \s_mux_signals[0][15][0] ,
         \s_mux_signals[0][16][31] , \s_mux_signals[0][16][30] ,
         \s_mux_signals[0][16][29] , \s_mux_signals[0][16][28] ,
         \s_mux_signals[0][16][27] , \s_mux_signals[0][16][26] ,
         \s_mux_signals[0][16][25] , \s_mux_signals[0][16][24] ,
         \s_mux_signals[0][16][23] , \s_mux_signals[0][16][22] ,
         \s_mux_signals[0][16][21] , \s_mux_signals[0][16][20] ,
         \s_mux_signals[0][16][19] , \s_mux_signals[0][16][18] ,
         \s_mux_signals[0][16][17] , \s_mux_signals[0][16][16] ,
         \s_mux_signals[0][16][15] , \s_mux_signals[0][16][14] ,
         \s_mux_signals[0][16][13] , \s_mux_signals[0][16][12] ,
         \s_mux_signals[0][16][11] , \s_mux_signals[0][16][10] ,
         \s_mux_signals[0][16][9] , \s_mux_signals[0][16][8] ,
         \s_mux_signals[0][16][7] , \s_mux_signals[0][16][6] ,
         \s_mux_signals[0][16][5] , \s_mux_signals[0][16][4] ,
         \s_mux_signals[0][16][3] , \s_mux_signals[0][16][2] ,
         \s_mux_signals[0][16][1] , \s_mux_signals[0][16][0] ,
         \s_mux_signals[0][17][31] , \s_mux_signals[0][17][30] ,
         \s_mux_signals[0][17][29] , \s_mux_signals[0][17][28] ,
         \s_mux_signals[0][17][27] , \s_mux_signals[0][17][26] ,
         \s_mux_signals[0][17][25] , \s_mux_signals[0][17][24] ,
         \s_mux_signals[0][17][23] , \s_mux_signals[0][17][22] ,
         \s_mux_signals[0][17][21] , \s_mux_signals[0][17][20] ,
         \s_mux_signals[0][17][19] , \s_mux_signals[0][17][18] ,
         \s_mux_signals[0][17][17] , \s_mux_signals[0][17][16] ,
         \s_mux_signals[0][17][15] , \s_mux_signals[0][17][14] ,
         \s_mux_signals[0][17][13] , \s_mux_signals[0][17][12] ,
         \s_mux_signals[0][17][11] , \s_mux_signals[0][17][10] ,
         \s_mux_signals[0][17][9] , \s_mux_signals[0][17][8] ,
         \s_mux_signals[0][17][7] , \s_mux_signals[0][17][6] ,
         \s_mux_signals[0][17][5] , \s_mux_signals[0][17][4] ,
         \s_mux_signals[0][17][3] , \s_mux_signals[0][17][2] ,
         \s_mux_signals[0][17][1] , \s_mux_signals[0][17][0] ,
         \s_mux_signals[0][18][31] , \s_mux_signals[0][18][30] ,
         \s_mux_signals[0][18][29] , \s_mux_signals[0][18][28] ,
         \s_mux_signals[0][18][27] , \s_mux_signals[0][18][26] ,
         \s_mux_signals[0][18][25] , \s_mux_signals[0][18][24] ,
         \s_mux_signals[0][18][23] , \s_mux_signals[0][18][22] ,
         \s_mux_signals[0][18][21] , \s_mux_signals[0][18][20] ,
         \s_mux_signals[0][18][19] , \s_mux_signals[0][18][18] ,
         \s_mux_signals[0][18][17] , \s_mux_signals[0][18][16] ,
         \s_mux_signals[0][18][15] , \s_mux_signals[0][18][14] ,
         \s_mux_signals[0][18][13] , \s_mux_signals[0][18][12] ,
         \s_mux_signals[0][18][11] , \s_mux_signals[0][18][10] ,
         \s_mux_signals[0][18][9] , \s_mux_signals[0][18][8] ,
         \s_mux_signals[0][18][7] , \s_mux_signals[0][18][6] ,
         \s_mux_signals[0][18][5] , \s_mux_signals[0][18][4] ,
         \s_mux_signals[0][18][3] , \s_mux_signals[0][18][2] ,
         \s_mux_signals[0][18][1] , \s_mux_signals[0][18][0] ,
         \s_mux_signals[0][19][31] , \s_mux_signals[0][19][30] ,
         \s_mux_signals[0][19][29] , \s_mux_signals[0][19][28] ,
         \s_mux_signals[0][19][27] , \s_mux_signals[0][19][26] ,
         \s_mux_signals[0][19][25] , \s_mux_signals[0][19][24] ,
         \s_mux_signals[0][19][23] , \s_mux_signals[0][19][22] ,
         \s_mux_signals[0][19][21] , \s_mux_signals[0][19][20] ,
         \s_mux_signals[0][19][19] , \s_mux_signals[0][19][18] ,
         \s_mux_signals[0][19][17] , \s_mux_signals[0][19][16] ,
         \s_mux_signals[0][19][15] , \s_mux_signals[0][19][14] ,
         \s_mux_signals[0][19][13] , \s_mux_signals[0][19][12] ,
         \s_mux_signals[0][19][11] , \s_mux_signals[0][19][10] ,
         \s_mux_signals[0][19][9] , \s_mux_signals[0][19][8] ,
         \s_mux_signals[0][19][7] , \s_mux_signals[0][19][6] ,
         \s_mux_signals[0][19][5] , \s_mux_signals[0][19][4] ,
         \s_mux_signals[0][19][3] , \s_mux_signals[0][19][2] ,
         \s_mux_signals[0][19][1] , \s_mux_signals[0][19][0] ,
         \s_mux_signals[0][20][31] , \s_mux_signals[0][20][30] ,
         \s_mux_signals[0][20][29] , \s_mux_signals[0][20][28] ,
         \s_mux_signals[0][20][27] , \s_mux_signals[0][20][26] ,
         \s_mux_signals[0][20][25] , \s_mux_signals[0][20][24] ,
         \s_mux_signals[0][20][23] , \s_mux_signals[0][20][22] ,
         \s_mux_signals[0][20][21] , \s_mux_signals[0][20][20] ,
         \s_mux_signals[0][20][19] , \s_mux_signals[0][20][18] ,
         \s_mux_signals[0][20][17] , \s_mux_signals[0][20][16] ,
         \s_mux_signals[0][20][15] , \s_mux_signals[0][20][14] ,
         \s_mux_signals[0][20][13] , \s_mux_signals[0][20][12] ,
         \s_mux_signals[0][20][11] , \s_mux_signals[0][20][10] ,
         \s_mux_signals[0][20][9] , \s_mux_signals[0][20][8] ,
         \s_mux_signals[0][20][7] , \s_mux_signals[0][20][6] ,
         \s_mux_signals[0][20][5] , \s_mux_signals[0][20][4] ,
         \s_mux_signals[0][20][3] , \s_mux_signals[0][20][2] ,
         \s_mux_signals[0][20][1] , \s_mux_signals[0][20][0] ,
         \s_mux_signals[0][21][31] , \s_mux_signals[0][21][30] ,
         \s_mux_signals[0][21][29] , \s_mux_signals[0][21][28] ,
         \s_mux_signals[0][21][27] , \s_mux_signals[0][21][26] ,
         \s_mux_signals[0][21][25] , \s_mux_signals[0][21][24] ,
         \s_mux_signals[0][21][23] , \s_mux_signals[0][21][22] ,
         \s_mux_signals[0][21][21] , \s_mux_signals[0][21][20] ,
         \s_mux_signals[0][21][19] , \s_mux_signals[0][21][18] ,
         \s_mux_signals[0][21][17] , \s_mux_signals[0][21][16] ,
         \s_mux_signals[0][21][15] , \s_mux_signals[0][21][14] ,
         \s_mux_signals[0][21][13] , \s_mux_signals[0][21][12] ,
         \s_mux_signals[0][21][11] , \s_mux_signals[0][21][10] ,
         \s_mux_signals[0][21][9] , \s_mux_signals[0][21][8] ,
         \s_mux_signals[0][21][7] , \s_mux_signals[0][21][6] ,
         \s_mux_signals[0][21][5] , \s_mux_signals[0][21][4] ,
         \s_mux_signals[0][21][3] , \s_mux_signals[0][21][2] ,
         \s_mux_signals[0][21][1] , \s_mux_signals[0][21][0] ,
         \s_mux_signals[0][22][31] , \s_mux_signals[0][22][30] ,
         \s_mux_signals[0][22][29] , \s_mux_signals[0][22][28] ,
         \s_mux_signals[0][22][27] , \s_mux_signals[0][22][26] ,
         \s_mux_signals[0][22][25] , \s_mux_signals[0][22][24] ,
         \s_mux_signals[0][22][23] , \s_mux_signals[0][22][22] ,
         \s_mux_signals[0][22][21] , \s_mux_signals[0][22][20] ,
         \s_mux_signals[0][22][19] , \s_mux_signals[0][22][18] ,
         \s_mux_signals[0][22][17] , \s_mux_signals[0][22][16] ,
         \s_mux_signals[0][22][15] , \s_mux_signals[0][22][14] ,
         \s_mux_signals[0][22][13] , \s_mux_signals[0][22][12] ,
         \s_mux_signals[0][22][11] , \s_mux_signals[0][22][10] ,
         \s_mux_signals[0][22][9] , \s_mux_signals[0][22][8] ,
         \s_mux_signals[0][22][7] , \s_mux_signals[0][22][6] ,
         \s_mux_signals[0][22][5] , \s_mux_signals[0][22][4] ,
         \s_mux_signals[0][22][3] , \s_mux_signals[0][22][2] ,
         \s_mux_signals[0][22][1] , \s_mux_signals[0][22][0] ,
         \s_mux_signals[0][23][31] , \s_mux_signals[0][23][30] ,
         \s_mux_signals[0][23][29] , \s_mux_signals[0][23][28] ,
         \s_mux_signals[0][23][27] , \s_mux_signals[0][23][26] ,
         \s_mux_signals[0][23][25] , \s_mux_signals[0][23][24] ,
         \s_mux_signals[0][23][23] , \s_mux_signals[0][23][22] ,
         \s_mux_signals[0][23][21] , \s_mux_signals[0][23][20] ,
         \s_mux_signals[0][23][19] , \s_mux_signals[0][23][18] ,
         \s_mux_signals[0][23][17] , \s_mux_signals[0][23][16] ,
         \s_mux_signals[0][23][15] , \s_mux_signals[0][23][14] ,
         \s_mux_signals[0][23][13] , \s_mux_signals[0][23][12] ,
         \s_mux_signals[0][23][11] , \s_mux_signals[0][23][10] ,
         \s_mux_signals[0][23][9] , \s_mux_signals[0][23][8] ,
         \s_mux_signals[0][23][7] , \s_mux_signals[0][23][6] ,
         \s_mux_signals[0][23][5] , \s_mux_signals[0][23][4] ,
         \s_mux_signals[0][23][3] , \s_mux_signals[0][23][2] ,
         \s_mux_signals[0][23][1] , \s_mux_signals[0][23][0] ,
         \s_mux_signals[0][24][31] , \s_mux_signals[0][24][30] ,
         \s_mux_signals[0][24][29] , \s_mux_signals[0][24][28] ,
         \s_mux_signals[0][24][27] , \s_mux_signals[0][24][26] ,
         \s_mux_signals[0][24][25] , \s_mux_signals[0][24][24] ,
         \s_mux_signals[0][24][23] , \s_mux_signals[0][24][22] ,
         \s_mux_signals[0][24][21] , \s_mux_signals[0][24][20] ,
         \s_mux_signals[0][24][19] , \s_mux_signals[0][24][18] ,
         \s_mux_signals[0][24][17] , \s_mux_signals[0][24][16] ,
         \s_mux_signals[0][24][15] , \s_mux_signals[0][24][14] ,
         \s_mux_signals[0][24][13] , \s_mux_signals[0][24][12] ,
         \s_mux_signals[0][24][11] , \s_mux_signals[0][24][10] ,
         \s_mux_signals[0][24][9] , \s_mux_signals[0][24][8] ,
         \s_mux_signals[0][24][7] , \s_mux_signals[0][24][6] ,
         \s_mux_signals[0][24][5] , \s_mux_signals[0][24][4] ,
         \s_mux_signals[0][24][3] , \s_mux_signals[0][24][2] ,
         \s_mux_signals[0][24][1] , \s_mux_signals[0][24][0] ,
         \s_mux_signals[0][25][31] , \s_mux_signals[0][25][30] ,
         \s_mux_signals[0][25][29] , \s_mux_signals[0][25][28] ,
         \s_mux_signals[0][25][27] , \s_mux_signals[0][25][26] ,
         \s_mux_signals[0][25][25] , \s_mux_signals[0][25][24] ,
         \s_mux_signals[0][25][23] , \s_mux_signals[0][25][22] ,
         \s_mux_signals[0][25][21] , \s_mux_signals[0][25][20] ,
         \s_mux_signals[0][25][19] , \s_mux_signals[0][25][18] ,
         \s_mux_signals[0][25][17] , \s_mux_signals[0][25][16] ,
         \s_mux_signals[0][25][15] , \s_mux_signals[0][25][14] ,
         \s_mux_signals[0][25][13] , \s_mux_signals[0][25][12] ,
         \s_mux_signals[0][25][11] , \s_mux_signals[0][25][10] ,
         \s_mux_signals[0][25][9] , \s_mux_signals[0][25][8] ,
         \s_mux_signals[0][25][7] , \s_mux_signals[0][25][6] ,
         \s_mux_signals[0][25][5] , \s_mux_signals[0][25][4] ,
         \s_mux_signals[0][25][3] , \s_mux_signals[0][25][2] ,
         \s_mux_signals[0][25][1] , \s_mux_signals[0][25][0] ,
         \s_mux_signals[0][26][31] , \s_mux_signals[0][26][30] ,
         \s_mux_signals[0][26][29] , \s_mux_signals[0][26][28] ,
         \s_mux_signals[0][26][27] , \s_mux_signals[0][26][26] ,
         \s_mux_signals[0][26][25] , \s_mux_signals[0][26][24] ,
         \s_mux_signals[0][26][23] , \s_mux_signals[0][26][22] ,
         \s_mux_signals[0][26][21] , \s_mux_signals[0][26][20] ,
         \s_mux_signals[0][26][19] , \s_mux_signals[0][26][18] ,
         \s_mux_signals[0][26][17] , \s_mux_signals[0][26][16] ,
         \s_mux_signals[0][26][15] , \s_mux_signals[0][26][14] ,
         \s_mux_signals[0][26][13] , \s_mux_signals[0][26][12] ,
         \s_mux_signals[0][26][11] , \s_mux_signals[0][26][10] ,
         \s_mux_signals[0][26][9] , \s_mux_signals[0][26][8] ,
         \s_mux_signals[0][26][7] , \s_mux_signals[0][26][6] ,
         \s_mux_signals[0][26][5] , \s_mux_signals[0][26][4] ,
         \s_mux_signals[0][26][3] , \s_mux_signals[0][26][2] ,
         \s_mux_signals[0][26][1] , \s_mux_signals[0][26][0] ,
         \s_mux_signals[0][27][31] , \s_mux_signals[0][27][30] ,
         \s_mux_signals[0][27][29] , \s_mux_signals[0][27][28] ,
         \s_mux_signals[0][27][27] , \s_mux_signals[0][27][26] ,
         \s_mux_signals[0][27][25] , \s_mux_signals[0][27][24] ,
         \s_mux_signals[0][27][23] , \s_mux_signals[0][27][22] ,
         \s_mux_signals[0][27][21] , \s_mux_signals[0][27][20] ,
         \s_mux_signals[0][27][19] , \s_mux_signals[0][27][18] ,
         \s_mux_signals[0][27][17] , \s_mux_signals[0][27][16] ,
         \s_mux_signals[0][27][15] , \s_mux_signals[0][27][14] ,
         \s_mux_signals[0][27][13] , \s_mux_signals[0][27][12] ,
         \s_mux_signals[0][27][11] , \s_mux_signals[0][27][10] ,
         \s_mux_signals[0][27][9] , \s_mux_signals[0][27][8] ,
         \s_mux_signals[0][27][7] , \s_mux_signals[0][27][6] ,
         \s_mux_signals[0][27][5] , \s_mux_signals[0][27][4] ,
         \s_mux_signals[0][27][3] , \s_mux_signals[0][27][2] ,
         \s_mux_signals[0][27][1] , \s_mux_signals[0][27][0] ,
         \s_mux_signals[0][28][31] , \s_mux_signals[0][28][30] ,
         \s_mux_signals[0][28][29] , \s_mux_signals[0][28][28] ,
         \s_mux_signals[0][28][27] , \s_mux_signals[0][28][26] ,
         \s_mux_signals[0][28][25] , \s_mux_signals[0][28][24] ,
         \s_mux_signals[0][28][23] , \s_mux_signals[0][28][22] ,
         \s_mux_signals[0][28][21] , \s_mux_signals[0][28][20] ,
         \s_mux_signals[0][28][19] , \s_mux_signals[0][28][18] ,
         \s_mux_signals[0][28][17] , \s_mux_signals[0][28][16] ,
         \s_mux_signals[0][28][15] , \s_mux_signals[0][28][14] ,
         \s_mux_signals[0][28][13] , \s_mux_signals[0][28][12] ,
         \s_mux_signals[0][28][11] , \s_mux_signals[0][28][10] ,
         \s_mux_signals[0][28][9] , \s_mux_signals[0][28][8] ,
         \s_mux_signals[0][28][7] , \s_mux_signals[0][28][6] ,
         \s_mux_signals[0][28][5] , \s_mux_signals[0][28][4] ,
         \s_mux_signals[0][28][3] , \s_mux_signals[0][28][2] ,
         \s_mux_signals[0][28][1] , \s_mux_signals[0][28][0] ,
         \s_mux_signals[0][29][31] , \s_mux_signals[0][29][30] ,
         \s_mux_signals[0][29][29] , \s_mux_signals[0][29][28] ,
         \s_mux_signals[0][29][27] , \s_mux_signals[0][29][26] ,
         \s_mux_signals[0][29][25] , \s_mux_signals[0][29][24] ,
         \s_mux_signals[0][29][23] , \s_mux_signals[0][29][22] ,
         \s_mux_signals[0][29][21] , \s_mux_signals[0][29][20] ,
         \s_mux_signals[0][29][19] , \s_mux_signals[0][29][18] ,
         \s_mux_signals[0][29][17] , \s_mux_signals[0][29][16] ,
         \s_mux_signals[0][29][15] , \s_mux_signals[0][29][14] ,
         \s_mux_signals[0][29][13] , \s_mux_signals[0][29][12] ,
         \s_mux_signals[0][29][11] , \s_mux_signals[0][29][10] ,
         \s_mux_signals[0][29][9] , \s_mux_signals[0][29][8] ,
         \s_mux_signals[0][29][7] , \s_mux_signals[0][29][6] ,
         \s_mux_signals[0][29][5] , \s_mux_signals[0][29][4] ,
         \s_mux_signals[0][29][3] , \s_mux_signals[0][29][2] ,
         \s_mux_signals[0][29][1] , \s_mux_signals[0][29][0] ,
         \s_mux_signals[0][30][31] , \s_mux_signals[0][30][30] ,
         \s_mux_signals[0][30][29] , \s_mux_signals[0][30][28] ,
         \s_mux_signals[0][30][27] , \s_mux_signals[0][30][26] ,
         \s_mux_signals[0][30][25] , \s_mux_signals[0][30][24] ,
         \s_mux_signals[0][30][23] , \s_mux_signals[0][30][22] ,
         \s_mux_signals[0][30][21] , \s_mux_signals[0][30][20] ,
         \s_mux_signals[0][30][19] , \s_mux_signals[0][30][18] ,
         \s_mux_signals[0][30][17] , \s_mux_signals[0][30][16] ,
         \s_mux_signals[0][30][15] , \s_mux_signals[0][30][14] ,
         \s_mux_signals[0][30][13] , \s_mux_signals[0][30][12] ,
         \s_mux_signals[0][30][11] , \s_mux_signals[0][30][10] ,
         \s_mux_signals[0][30][9] , \s_mux_signals[0][30][8] ,
         \s_mux_signals[0][30][7] , \s_mux_signals[0][30][6] ,
         \s_mux_signals[0][30][5] , \s_mux_signals[0][30][4] ,
         \s_mux_signals[0][30][3] , \s_mux_signals[0][30][2] ,
         \s_mux_signals[0][30][1] , \s_mux_signals[0][30][0] ,
         \s_mux_signals[0][31][31] , \s_mux_signals[0][31][30] ,
         \s_mux_signals[0][31][29] , \s_mux_signals[0][31][28] ,
         \s_mux_signals[0][31][27] , \s_mux_signals[0][31][26] ,
         \s_mux_signals[0][31][25] , \s_mux_signals[0][31][24] ,
         \s_mux_signals[0][31][23] , \s_mux_signals[0][31][22] ,
         \s_mux_signals[0][31][21] , \s_mux_signals[0][31][20] ,
         \s_mux_signals[0][31][19] , \s_mux_signals[0][31][18] ,
         \s_mux_signals[0][31][17] , \s_mux_signals[0][31][16] ,
         \s_mux_signals[0][31][15] , \s_mux_signals[0][31][14] ,
         \s_mux_signals[0][31][13] , \s_mux_signals[0][31][12] ,
         \s_mux_signals[0][31][11] , \s_mux_signals[0][31][10] ,
         \s_mux_signals[0][31][9] , \s_mux_signals[0][31][8] ,
         \s_mux_signals[0][31][7] , \s_mux_signals[0][31][6] ,
         \s_mux_signals[0][31][5] , \s_mux_signals[0][31][4] ,
         \s_mux_signals[0][31][3] , \s_mux_signals[0][31][2] ,
         \s_mux_signals[0][31][1] , \s_mux_signals[0][31][0] ,
         \s_mux_signals[1][0][31] , \s_mux_signals[1][0][30] ,
         \s_mux_signals[1][0][29] , \s_mux_signals[1][0][28] ,
         \s_mux_signals[1][0][27] , \s_mux_signals[1][0][26] ,
         \s_mux_signals[1][0][25] , \s_mux_signals[1][0][24] ,
         \s_mux_signals[1][0][23] , \s_mux_signals[1][0][22] ,
         \s_mux_signals[1][0][21] , \s_mux_signals[1][0][20] ,
         \s_mux_signals[1][0][19] , \s_mux_signals[1][0][18] ,
         \s_mux_signals[1][0][17] , \s_mux_signals[1][0][16] ,
         \s_mux_signals[1][0][15] , \s_mux_signals[1][0][14] ,
         \s_mux_signals[1][0][13] , \s_mux_signals[1][0][12] ,
         \s_mux_signals[1][0][11] , \s_mux_signals[1][0][10] ,
         \s_mux_signals[1][0][9] , \s_mux_signals[1][0][8] ,
         \s_mux_signals[1][0][7] , \s_mux_signals[1][0][6] ,
         \s_mux_signals[1][0][5] , \s_mux_signals[1][0][4] ,
         \s_mux_signals[1][0][3] , \s_mux_signals[1][0][2] ,
         \s_mux_signals[1][0][1] , \s_mux_signals[1][0][0] ,
         \s_mux_signals[1][2][31] , \s_mux_signals[1][2][30] ,
         \s_mux_signals[1][2][29] , \s_mux_signals[1][2][28] ,
         \s_mux_signals[1][2][27] , \s_mux_signals[1][2][26] ,
         \s_mux_signals[1][2][25] , \s_mux_signals[1][2][24] ,
         \s_mux_signals[1][2][23] , \s_mux_signals[1][2][22] ,
         \s_mux_signals[1][2][21] , \s_mux_signals[1][2][20] ,
         \s_mux_signals[1][2][19] , \s_mux_signals[1][2][18] ,
         \s_mux_signals[1][2][17] , \s_mux_signals[1][2][16] ,
         \s_mux_signals[1][2][15] , \s_mux_signals[1][2][14] ,
         \s_mux_signals[1][2][13] , \s_mux_signals[1][2][12] ,
         \s_mux_signals[1][2][11] , \s_mux_signals[1][2][10] ,
         \s_mux_signals[1][2][9] , \s_mux_signals[1][2][8] ,
         \s_mux_signals[1][2][7] , \s_mux_signals[1][2][6] ,
         \s_mux_signals[1][2][5] , \s_mux_signals[1][2][4] ,
         \s_mux_signals[1][2][3] , \s_mux_signals[1][2][2] ,
         \s_mux_signals[1][2][1] , \s_mux_signals[1][2][0] ,
         \s_mux_signals[1][4][31] , \s_mux_signals[1][4][30] ,
         \s_mux_signals[1][4][29] , \s_mux_signals[1][4][28] ,
         \s_mux_signals[1][4][27] , \s_mux_signals[1][4][26] ,
         \s_mux_signals[1][4][25] , \s_mux_signals[1][4][24] ,
         \s_mux_signals[1][4][23] , \s_mux_signals[1][4][22] ,
         \s_mux_signals[1][4][21] , \s_mux_signals[1][4][20] ,
         \s_mux_signals[1][4][19] , \s_mux_signals[1][4][18] ,
         \s_mux_signals[1][4][17] , \s_mux_signals[1][4][16] ,
         \s_mux_signals[1][4][15] , \s_mux_signals[1][4][14] ,
         \s_mux_signals[1][4][13] , \s_mux_signals[1][4][12] ,
         \s_mux_signals[1][4][11] , \s_mux_signals[1][4][10] ,
         \s_mux_signals[1][4][9] , \s_mux_signals[1][4][8] ,
         \s_mux_signals[1][4][7] , \s_mux_signals[1][4][6] ,
         \s_mux_signals[1][4][5] , \s_mux_signals[1][4][4] ,
         \s_mux_signals[1][4][3] , \s_mux_signals[1][4][2] ,
         \s_mux_signals[1][4][1] , \s_mux_signals[1][4][0] ,
         \s_mux_signals[1][6][31] , \s_mux_signals[1][6][30] ,
         \s_mux_signals[1][6][29] , \s_mux_signals[1][6][28] ,
         \s_mux_signals[1][6][27] , \s_mux_signals[1][6][26] ,
         \s_mux_signals[1][6][25] , \s_mux_signals[1][6][24] ,
         \s_mux_signals[1][6][23] , \s_mux_signals[1][6][22] ,
         \s_mux_signals[1][6][21] , \s_mux_signals[1][6][20] ,
         \s_mux_signals[1][6][19] , \s_mux_signals[1][6][18] ,
         \s_mux_signals[1][6][17] , \s_mux_signals[1][6][16] ,
         \s_mux_signals[1][6][15] , \s_mux_signals[1][6][14] ,
         \s_mux_signals[1][6][13] , \s_mux_signals[1][6][12] ,
         \s_mux_signals[1][6][11] , \s_mux_signals[1][6][10] ,
         \s_mux_signals[1][6][9] , \s_mux_signals[1][6][8] ,
         \s_mux_signals[1][6][7] , \s_mux_signals[1][6][6] ,
         \s_mux_signals[1][6][5] , \s_mux_signals[1][6][4] ,
         \s_mux_signals[1][6][3] , \s_mux_signals[1][6][2] ,
         \s_mux_signals[1][6][1] , \s_mux_signals[1][6][0] ,
         \s_mux_signals[1][8][31] , \s_mux_signals[1][8][30] ,
         \s_mux_signals[1][8][29] , \s_mux_signals[1][8][28] ,
         \s_mux_signals[1][8][27] , \s_mux_signals[1][8][26] ,
         \s_mux_signals[1][8][25] , \s_mux_signals[1][8][24] ,
         \s_mux_signals[1][8][23] , \s_mux_signals[1][8][22] ,
         \s_mux_signals[1][8][21] , \s_mux_signals[1][8][20] ,
         \s_mux_signals[1][8][19] , \s_mux_signals[1][8][18] ,
         \s_mux_signals[1][8][17] , \s_mux_signals[1][8][16] ,
         \s_mux_signals[1][8][15] , \s_mux_signals[1][8][14] ,
         \s_mux_signals[1][8][13] , \s_mux_signals[1][8][12] ,
         \s_mux_signals[1][8][11] , \s_mux_signals[1][8][10] ,
         \s_mux_signals[1][8][9] , \s_mux_signals[1][8][8] ,
         \s_mux_signals[1][8][7] , \s_mux_signals[1][8][6] ,
         \s_mux_signals[1][8][5] , \s_mux_signals[1][8][4] ,
         \s_mux_signals[1][8][3] , \s_mux_signals[1][8][2] ,
         \s_mux_signals[1][8][1] , \s_mux_signals[1][8][0] ,
         \s_mux_signals[1][10][31] , \s_mux_signals[1][10][30] ,
         \s_mux_signals[1][10][29] , \s_mux_signals[1][10][28] ,
         \s_mux_signals[1][10][27] , \s_mux_signals[1][10][26] ,
         \s_mux_signals[1][10][25] , \s_mux_signals[1][10][24] ,
         \s_mux_signals[1][10][23] , \s_mux_signals[1][10][22] ,
         \s_mux_signals[1][10][21] , \s_mux_signals[1][10][20] ,
         \s_mux_signals[1][10][19] , \s_mux_signals[1][10][18] ,
         \s_mux_signals[1][10][17] , \s_mux_signals[1][10][16] ,
         \s_mux_signals[1][10][15] , \s_mux_signals[1][10][14] ,
         \s_mux_signals[1][10][13] , \s_mux_signals[1][10][12] ,
         \s_mux_signals[1][10][11] , \s_mux_signals[1][10][10] ,
         \s_mux_signals[1][10][9] , \s_mux_signals[1][10][8] ,
         \s_mux_signals[1][10][7] , \s_mux_signals[1][10][6] ,
         \s_mux_signals[1][10][5] , \s_mux_signals[1][10][4] ,
         \s_mux_signals[1][10][3] , \s_mux_signals[1][10][2] ,
         \s_mux_signals[1][10][1] , \s_mux_signals[1][10][0] ,
         \s_mux_signals[1][12][31] , \s_mux_signals[1][12][30] ,
         \s_mux_signals[1][12][29] , \s_mux_signals[1][12][28] ,
         \s_mux_signals[1][12][27] , \s_mux_signals[1][12][26] ,
         \s_mux_signals[1][12][25] , \s_mux_signals[1][12][24] ,
         \s_mux_signals[1][12][23] , \s_mux_signals[1][12][22] ,
         \s_mux_signals[1][12][21] , \s_mux_signals[1][12][20] ,
         \s_mux_signals[1][12][19] , \s_mux_signals[1][12][18] ,
         \s_mux_signals[1][12][17] , \s_mux_signals[1][12][16] ,
         \s_mux_signals[1][12][15] , \s_mux_signals[1][12][14] ,
         \s_mux_signals[1][12][13] , \s_mux_signals[1][12][12] ,
         \s_mux_signals[1][12][11] , \s_mux_signals[1][12][10] ,
         \s_mux_signals[1][12][9] , \s_mux_signals[1][12][8] ,
         \s_mux_signals[1][12][7] , \s_mux_signals[1][12][6] ,
         \s_mux_signals[1][12][5] , \s_mux_signals[1][12][4] ,
         \s_mux_signals[1][12][3] , \s_mux_signals[1][12][2] ,
         \s_mux_signals[1][12][1] , \s_mux_signals[1][12][0] ,
         \s_mux_signals[1][14][31] , \s_mux_signals[1][14][30] ,
         \s_mux_signals[1][14][29] , \s_mux_signals[1][14][28] ,
         \s_mux_signals[1][14][27] , \s_mux_signals[1][14][26] ,
         \s_mux_signals[1][14][25] , \s_mux_signals[1][14][24] ,
         \s_mux_signals[1][14][23] , \s_mux_signals[1][14][22] ,
         \s_mux_signals[1][14][21] , \s_mux_signals[1][14][20] ,
         \s_mux_signals[1][14][19] , \s_mux_signals[1][14][18] ,
         \s_mux_signals[1][14][17] , \s_mux_signals[1][14][16] ,
         \s_mux_signals[1][14][15] , \s_mux_signals[1][14][14] ,
         \s_mux_signals[1][14][13] , \s_mux_signals[1][14][12] ,
         \s_mux_signals[1][14][11] , \s_mux_signals[1][14][10] ,
         \s_mux_signals[1][14][9] , \s_mux_signals[1][14][8] ,
         \s_mux_signals[1][14][7] , \s_mux_signals[1][14][6] ,
         \s_mux_signals[1][14][5] , \s_mux_signals[1][14][4] ,
         \s_mux_signals[1][14][3] , \s_mux_signals[1][14][2] ,
         \s_mux_signals[1][14][1] , \s_mux_signals[1][14][0] ,
         \s_mux_signals[1][16][31] , \s_mux_signals[1][16][30] ,
         \s_mux_signals[1][16][29] , \s_mux_signals[1][16][28] ,
         \s_mux_signals[1][16][27] , \s_mux_signals[1][16][26] ,
         \s_mux_signals[1][16][25] , \s_mux_signals[1][16][24] ,
         \s_mux_signals[1][16][23] , \s_mux_signals[1][16][22] ,
         \s_mux_signals[1][16][21] , \s_mux_signals[1][16][20] ,
         \s_mux_signals[1][16][19] , \s_mux_signals[1][16][18] ,
         \s_mux_signals[1][16][17] , \s_mux_signals[1][16][16] ,
         \s_mux_signals[1][16][15] , \s_mux_signals[1][16][14] ,
         \s_mux_signals[1][16][13] , \s_mux_signals[1][16][12] ,
         \s_mux_signals[1][16][11] , \s_mux_signals[1][16][10] ,
         \s_mux_signals[1][16][9] , \s_mux_signals[1][16][8] ,
         \s_mux_signals[1][16][7] , \s_mux_signals[1][16][6] ,
         \s_mux_signals[1][16][5] , \s_mux_signals[1][16][4] ,
         \s_mux_signals[1][16][3] , \s_mux_signals[1][16][2] ,
         \s_mux_signals[1][16][1] , \s_mux_signals[1][16][0] ,
         \s_mux_signals[1][18][31] , \s_mux_signals[1][18][30] ,
         \s_mux_signals[1][18][29] , \s_mux_signals[1][18][28] ,
         \s_mux_signals[1][18][27] , \s_mux_signals[1][18][26] ,
         \s_mux_signals[1][18][25] , \s_mux_signals[1][18][24] ,
         \s_mux_signals[1][18][23] , \s_mux_signals[1][18][22] ,
         \s_mux_signals[1][18][21] , \s_mux_signals[1][18][20] ,
         \s_mux_signals[1][18][19] , \s_mux_signals[1][18][18] ,
         \s_mux_signals[1][18][17] , \s_mux_signals[1][18][16] ,
         \s_mux_signals[1][18][15] , \s_mux_signals[1][18][14] ,
         \s_mux_signals[1][18][13] , \s_mux_signals[1][18][12] ,
         \s_mux_signals[1][18][11] , \s_mux_signals[1][18][10] ,
         \s_mux_signals[1][18][9] , \s_mux_signals[1][18][8] ,
         \s_mux_signals[1][18][7] , \s_mux_signals[1][18][6] ,
         \s_mux_signals[1][18][5] , \s_mux_signals[1][18][4] ,
         \s_mux_signals[1][18][3] , \s_mux_signals[1][18][2] ,
         \s_mux_signals[1][18][1] , \s_mux_signals[1][18][0] ,
         \s_mux_signals[1][20][31] , \s_mux_signals[1][20][30] ,
         \s_mux_signals[1][20][29] , \s_mux_signals[1][20][28] ,
         \s_mux_signals[1][20][27] , \s_mux_signals[1][20][26] ,
         \s_mux_signals[1][20][25] , \s_mux_signals[1][20][24] ,
         \s_mux_signals[1][20][23] , \s_mux_signals[1][20][22] ,
         \s_mux_signals[1][20][21] , \s_mux_signals[1][20][20] ,
         \s_mux_signals[1][20][19] , \s_mux_signals[1][20][18] ,
         \s_mux_signals[1][20][17] , \s_mux_signals[1][20][16] ,
         \s_mux_signals[1][20][15] , \s_mux_signals[1][20][14] ,
         \s_mux_signals[1][20][13] , \s_mux_signals[1][20][12] ,
         \s_mux_signals[1][20][11] , \s_mux_signals[1][20][10] ,
         \s_mux_signals[1][20][9] , \s_mux_signals[1][20][8] ,
         \s_mux_signals[1][20][7] , \s_mux_signals[1][20][6] ,
         \s_mux_signals[1][20][5] , \s_mux_signals[1][20][4] ,
         \s_mux_signals[1][20][3] , \s_mux_signals[1][20][2] ,
         \s_mux_signals[1][20][1] , \s_mux_signals[1][20][0] ,
         \s_mux_signals[1][22][31] , \s_mux_signals[1][22][30] ,
         \s_mux_signals[1][22][29] , \s_mux_signals[1][22][28] ,
         \s_mux_signals[1][22][27] , \s_mux_signals[1][22][26] ,
         \s_mux_signals[1][22][25] , \s_mux_signals[1][22][24] ,
         \s_mux_signals[1][22][23] , \s_mux_signals[1][22][22] ,
         \s_mux_signals[1][22][21] , \s_mux_signals[1][22][20] ,
         \s_mux_signals[1][22][19] , \s_mux_signals[1][22][18] ,
         \s_mux_signals[1][22][17] , \s_mux_signals[1][22][16] ,
         \s_mux_signals[1][22][15] , \s_mux_signals[1][22][14] ,
         \s_mux_signals[1][22][13] , \s_mux_signals[1][22][12] ,
         \s_mux_signals[1][22][11] , \s_mux_signals[1][22][10] ,
         \s_mux_signals[1][22][9] , \s_mux_signals[1][22][8] ,
         \s_mux_signals[1][22][7] , \s_mux_signals[1][22][6] ,
         \s_mux_signals[1][22][5] , \s_mux_signals[1][22][4] ,
         \s_mux_signals[1][22][3] , \s_mux_signals[1][22][2] ,
         \s_mux_signals[1][22][1] , \s_mux_signals[1][22][0] ,
         \s_mux_signals[1][24][31] , \s_mux_signals[1][24][30] ,
         \s_mux_signals[1][24][29] , \s_mux_signals[1][24][28] ,
         \s_mux_signals[1][24][27] , \s_mux_signals[1][24][26] ,
         \s_mux_signals[1][24][25] , \s_mux_signals[1][24][24] ,
         \s_mux_signals[1][24][23] , \s_mux_signals[1][24][22] ,
         \s_mux_signals[1][24][21] , \s_mux_signals[1][24][20] ,
         \s_mux_signals[1][24][19] , \s_mux_signals[1][24][18] ,
         \s_mux_signals[1][24][17] , \s_mux_signals[1][24][16] ,
         \s_mux_signals[1][24][15] , \s_mux_signals[1][24][14] ,
         \s_mux_signals[1][24][13] , \s_mux_signals[1][24][12] ,
         \s_mux_signals[1][24][11] , \s_mux_signals[1][24][10] ,
         \s_mux_signals[1][24][9] , \s_mux_signals[1][24][8] ,
         \s_mux_signals[1][24][7] , \s_mux_signals[1][24][6] ,
         \s_mux_signals[1][24][5] , \s_mux_signals[1][24][4] ,
         \s_mux_signals[1][24][3] , \s_mux_signals[1][24][2] ,
         \s_mux_signals[1][24][1] , \s_mux_signals[1][24][0] ,
         \s_mux_signals[1][26][31] , \s_mux_signals[1][26][30] ,
         \s_mux_signals[1][26][29] , \s_mux_signals[1][26][28] ,
         \s_mux_signals[1][26][27] , \s_mux_signals[1][26][26] ,
         \s_mux_signals[1][26][25] , \s_mux_signals[1][26][24] ,
         \s_mux_signals[1][26][23] , \s_mux_signals[1][26][22] ,
         \s_mux_signals[1][26][21] , \s_mux_signals[1][26][20] ,
         \s_mux_signals[1][26][19] , \s_mux_signals[1][26][18] ,
         \s_mux_signals[1][26][17] , \s_mux_signals[1][26][16] ,
         \s_mux_signals[1][26][15] , \s_mux_signals[1][26][14] ,
         \s_mux_signals[1][26][13] , \s_mux_signals[1][26][12] ,
         \s_mux_signals[1][26][11] , \s_mux_signals[1][26][10] ,
         \s_mux_signals[1][26][9] , \s_mux_signals[1][26][8] ,
         \s_mux_signals[1][26][7] , \s_mux_signals[1][26][6] ,
         \s_mux_signals[1][26][5] , \s_mux_signals[1][26][4] ,
         \s_mux_signals[1][26][3] , \s_mux_signals[1][26][2] ,
         \s_mux_signals[1][26][1] , \s_mux_signals[1][26][0] ,
         \s_mux_signals[1][28][31] , \s_mux_signals[1][28][30] ,
         \s_mux_signals[1][28][29] , \s_mux_signals[1][28][28] ,
         \s_mux_signals[1][28][27] , \s_mux_signals[1][28][26] ,
         \s_mux_signals[1][28][25] , \s_mux_signals[1][28][24] ,
         \s_mux_signals[1][28][23] , \s_mux_signals[1][28][22] ,
         \s_mux_signals[1][28][21] , \s_mux_signals[1][28][20] ,
         \s_mux_signals[1][28][19] , \s_mux_signals[1][28][18] ,
         \s_mux_signals[1][28][17] , \s_mux_signals[1][28][16] ,
         \s_mux_signals[1][28][15] , \s_mux_signals[1][28][14] ,
         \s_mux_signals[1][28][13] , \s_mux_signals[1][28][12] ,
         \s_mux_signals[1][28][11] , \s_mux_signals[1][28][10] ,
         \s_mux_signals[1][28][9] , \s_mux_signals[1][28][8] ,
         \s_mux_signals[1][28][7] , \s_mux_signals[1][28][6] ,
         \s_mux_signals[1][28][5] , \s_mux_signals[1][28][4] ,
         \s_mux_signals[1][28][3] , \s_mux_signals[1][28][2] ,
         \s_mux_signals[1][28][1] , \s_mux_signals[1][28][0] ,
         \s_mux_signals[1][30][31] , \s_mux_signals[1][30][30] ,
         \s_mux_signals[1][30][29] , \s_mux_signals[1][30][28] ,
         \s_mux_signals[1][30][27] , \s_mux_signals[1][30][26] ,
         \s_mux_signals[1][30][25] , \s_mux_signals[1][30][24] ,
         \s_mux_signals[1][30][23] , \s_mux_signals[1][30][22] ,
         \s_mux_signals[1][30][21] , \s_mux_signals[1][30][20] ,
         \s_mux_signals[1][30][19] , \s_mux_signals[1][30][18] ,
         \s_mux_signals[1][30][17] , \s_mux_signals[1][30][16] ,
         \s_mux_signals[1][30][15] , \s_mux_signals[1][30][14] ,
         \s_mux_signals[1][30][13] , \s_mux_signals[1][30][12] ,
         \s_mux_signals[1][30][11] , \s_mux_signals[1][30][10] ,
         \s_mux_signals[1][30][9] , \s_mux_signals[1][30][8] ,
         \s_mux_signals[1][30][7] , \s_mux_signals[1][30][6] ,
         \s_mux_signals[1][30][5] , \s_mux_signals[1][30][4] ,
         \s_mux_signals[1][30][3] , \s_mux_signals[1][30][2] ,
         \s_mux_signals[1][30][1] , \s_mux_signals[1][30][0] ,
         \s_mux_signals[2][0][31] , \s_mux_signals[2][0][30] ,
         \s_mux_signals[2][0][29] , \s_mux_signals[2][0][28] ,
         \s_mux_signals[2][0][27] , \s_mux_signals[2][0][26] ,
         \s_mux_signals[2][0][25] , \s_mux_signals[2][0][24] ,
         \s_mux_signals[2][0][23] , \s_mux_signals[2][0][22] ,
         \s_mux_signals[2][0][21] , \s_mux_signals[2][0][20] ,
         \s_mux_signals[2][0][19] , \s_mux_signals[2][0][18] ,
         \s_mux_signals[2][0][17] , \s_mux_signals[2][0][16] ,
         \s_mux_signals[2][0][15] , \s_mux_signals[2][0][14] ,
         \s_mux_signals[2][0][13] , \s_mux_signals[2][0][12] ,
         \s_mux_signals[2][0][11] , \s_mux_signals[2][0][10] ,
         \s_mux_signals[2][0][9] , \s_mux_signals[2][0][8] ,
         \s_mux_signals[2][0][7] , \s_mux_signals[2][0][6] ,
         \s_mux_signals[2][0][5] , \s_mux_signals[2][0][4] ,
         \s_mux_signals[2][0][3] , \s_mux_signals[2][0][2] ,
         \s_mux_signals[2][0][1] , \s_mux_signals[2][0][0] ,
         \s_mux_signals[2][4][31] , \s_mux_signals[2][4][30] ,
         \s_mux_signals[2][4][29] , \s_mux_signals[2][4][28] ,
         \s_mux_signals[2][4][27] , \s_mux_signals[2][4][26] ,
         \s_mux_signals[2][4][25] , \s_mux_signals[2][4][24] ,
         \s_mux_signals[2][4][23] , \s_mux_signals[2][4][22] ,
         \s_mux_signals[2][4][21] , \s_mux_signals[2][4][20] ,
         \s_mux_signals[2][4][19] , \s_mux_signals[2][4][18] ,
         \s_mux_signals[2][4][17] , \s_mux_signals[2][4][16] ,
         \s_mux_signals[2][4][15] , \s_mux_signals[2][4][14] ,
         \s_mux_signals[2][4][13] , \s_mux_signals[2][4][12] ,
         \s_mux_signals[2][4][11] , \s_mux_signals[2][4][10] ,
         \s_mux_signals[2][4][9] , \s_mux_signals[2][4][8] ,
         \s_mux_signals[2][4][7] , \s_mux_signals[2][4][6] ,
         \s_mux_signals[2][4][5] , \s_mux_signals[2][4][4] ,
         \s_mux_signals[2][4][3] , \s_mux_signals[2][4][2] ,
         \s_mux_signals[2][4][1] , \s_mux_signals[2][4][0] ,
         \s_mux_signals[2][8][31] , \s_mux_signals[2][8][30] ,
         \s_mux_signals[2][8][29] , \s_mux_signals[2][8][28] ,
         \s_mux_signals[2][8][27] , \s_mux_signals[2][8][26] ,
         \s_mux_signals[2][8][25] , \s_mux_signals[2][8][24] ,
         \s_mux_signals[2][8][23] , \s_mux_signals[2][8][22] ,
         \s_mux_signals[2][8][21] , \s_mux_signals[2][8][20] ,
         \s_mux_signals[2][8][19] , \s_mux_signals[2][8][18] ,
         \s_mux_signals[2][8][17] , \s_mux_signals[2][8][16] ,
         \s_mux_signals[2][8][15] , \s_mux_signals[2][8][14] ,
         \s_mux_signals[2][8][13] , \s_mux_signals[2][8][12] ,
         \s_mux_signals[2][8][11] , \s_mux_signals[2][8][10] ,
         \s_mux_signals[2][8][9] , \s_mux_signals[2][8][8] ,
         \s_mux_signals[2][8][7] , \s_mux_signals[2][8][6] ,
         \s_mux_signals[2][8][5] , \s_mux_signals[2][8][4] ,
         \s_mux_signals[2][8][3] , \s_mux_signals[2][8][2] ,
         \s_mux_signals[2][8][1] , \s_mux_signals[2][8][0] ,
         \s_mux_signals[2][12][31] , \s_mux_signals[2][12][30] ,
         \s_mux_signals[2][12][29] , \s_mux_signals[2][12][28] ,
         \s_mux_signals[2][12][27] , \s_mux_signals[2][12][26] ,
         \s_mux_signals[2][12][25] , \s_mux_signals[2][12][24] ,
         \s_mux_signals[2][12][23] , \s_mux_signals[2][12][22] ,
         \s_mux_signals[2][12][21] , \s_mux_signals[2][12][20] ,
         \s_mux_signals[2][12][19] , \s_mux_signals[2][12][18] ,
         \s_mux_signals[2][12][17] , \s_mux_signals[2][12][16] ,
         \s_mux_signals[2][12][15] , \s_mux_signals[2][12][14] ,
         \s_mux_signals[2][12][13] , \s_mux_signals[2][12][12] ,
         \s_mux_signals[2][12][11] , \s_mux_signals[2][12][10] ,
         \s_mux_signals[2][12][9] , \s_mux_signals[2][12][8] ,
         \s_mux_signals[2][12][7] , \s_mux_signals[2][12][6] ,
         \s_mux_signals[2][12][5] , \s_mux_signals[2][12][4] ,
         \s_mux_signals[2][12][3] , \s_mux_signals[2][12][2] ,
         \s_mux_signals[2][12][1] , \s_mux_signals[2][12][0] ,
         \s_mux_signals[2][16][31] , \s_mux_signals[2][16][30] ,
         \s_mux_signals[2][16][29] , \s_mux_signals[2][16][28] ,
         \s_mux_signals[2][16][27] , \s_mux_signals[2][16][26] ,
         \s_mux_signals[2][16][25] , \s_mux_signals[2][16][24] ,
         \s_mux_signals[2][16][23] , \s_mux_signals[2][16][22] ,
         \s_mux_signals[2][16][21] , \s_mux_signals[2][16][20] ,
         \s_mux_signals[2][16][19] , \s_mux_signals[2][16][18] ,
         \s_mux_signals[2][16][17] , \s_mux_signals[2][16][16] ,
         \s_mux_signals[2][16][15] , \s_mux_signals[2][16][14] ,
         \s_mux_signals[2][16][13] , \s_mux_signals[2][16][12] ,
         \s_mux_signals[2][16][11] , \s_mux_signals[2][16][10] ,
         \s_mux_signals[2][16][9] , \s_mux_signals[2][16][8] ,
         \s_mux_signals[2][16][7] , \s_mux_signals[2][16][6] ,
         \s_mux_signals[2][16][5] , \s_mux_signals[2][16][4] ,
         \s_mux_signals[2][16][3] , \s_mux_signals[2][16][2] ,
         \s_mux_signals[2][16][1] , \s_mux_signals[2][16][0] ,
         \s_mux_signals[2][20][31] , \s_mux_signals[2][20][30] ,
         \s_mux_signals[2][20][29] , \s_mux_signals[2][20][28] ,
         \s_mux_signals[2][20][27] , \s_mux_signals[2][20][26] ,
         \s_mux_signals[2][20][25] , \s_mux_signals[2][20][24] ,
         \s_mux_signals[2][20][23] , \s_mux_signals[2][20][22] ,
         \s_mux_signals[2][20][21] , \s_mux_signals[2][20][20] ,
         \s_mux_signals[2][20][19] , \s_mux_signals[2][20][18] ,
         \s_mux_signals[2][20][17] , \s_mux_signals[2][20][16] ,
         \s_mux_signals[2][20][15] , \s_mux_signals[2][20][14] ,
         \s_mux_signals[2][20][13] , \s_mux_signals[2][20][12] ,
         \s_mux_signals[2][20][11] , \s_mux_signals[2][20][10] ,
         \s_mux_signals[2][20][9] , \s_mux_signals[2][20][8] ,
         \s_mux_signals[2][20][7] , \s_mux_signals[2][20][6] ,
         \s_mux_signals[2][20][5] , \s_mux_signals[2][20][4] ,
         \s_mux_signals[2][20][3] , \s_mux_signals[2][20][2] ,
         \s_mux_signals[2][20][1] , \s_mux_signals[2][20][0] ,
         \s_mux_signals[2][24][31] , \s_mux_signals[2][24][30] ,
         \s_mux_signals[2][24][29] , \s_mux_signals[2][24][28] ,
         \s_mux_signals[2][24][27] , \s_mux_signals[2][24][26] ,
         \s_mux_signals[2][24][25] , \s_mux_signals[2][24][24] ,
         \s_mux_signals[2][24][23] , \s_mux_signals[2][24][22] ,
         \s_mux_signals[2][24][21] , \s_mux_signals[2][24][20] ,
         \s_mux_signals[2][24][19] , \s_mux_signals[2][24][18] ,
         \s_mux_signals[2][24][17] , \s_mux_signals[2][24][16] ,
         \s_mux_signals[2][24][15] , \s_mux_signals[2][24][14] ,
         \s_mux_signals[2][24][13] , \s_mux_signals[2][24][12] ,
         \s_mux_signals[2][24][11] , \s_mux_signals[2][24][10] ,
         \s_mux_signals[2][24][9] , \s_mux_signals[2][24][8] ,
         \s_mux_signals[2][24][7] , \s_mux_signals[2][24][6] ,
         \s_mux_signals[2][24][5] , \s_mux_signals[2][24][4] ,
         \s_mux_signals[2][24][3] , \s_mux_signals[2][24][2] ,
         \s_mux_signals[2][24][1] , \s_mux_signals[2][24][0] ,
         \s_mux_signals[2][28][31] , \s_mux_signals[2][28][30] ,
         \s_mux_signals[2][28][29] , \s_mux_signals[2][28][28] ,
         \s_mux_signals[2][28][27] , \s_mux_signals[2][28][26] ,
         \s_mux_signals[2][28][25] , \s_mux_signals[2][28][24] ,
         \s_mux_signals[2][28][23] , \s_mux_signals[2][28][22] ,
         \s_mux_signals[2][28][21] , \s_mux_signals[2][28][20] ,
         \s_mux_signals[2][28][19] , \s_mux_signals[2][28][18] ,
         \s_mux_signals[2][28][17] , \s_mux_signals[2][28][16] ,
         \s_mux_signals[2][28][15] , \s_mux_signals[2][28][14] ,
         \s_mux_signals[2][28][13] , \s_mux_signals[2][28][12] ,
         \s_mux_signals[2][28][11] , \s_mux_signals[2][28][10] ,
         \s_mux_signals[2][28][9] , \s_mux_signals[2][28][8] ,
         \s_mux_signals[2][28][7] , \s_mux_signals[2][28][6] ,
         \s_mux_signals[2][28][5] , \s_mux_signals[2][28][4] ,
         \s_mux_signals[2][28][3] , \s_mux_signals[2][28][2] ,
         \s_mux_signals[2][28][1] , \s_mux_signals[2][28][0] ,
         \s_mux_signals[3][0][31] , \s_mux_signals[3][0][30] ,
         \s_mux_signals[3][0][29] , \s_mux_signals[3][0][28] ,
         \s_mux_signals[3][0][27] , \s_mux_signals[3][0][26] ,
         \s_mux_signals[3][0][25] , \s_mux_signals[3][0][24] ,
         \s_mux_signals[3][0][23] , \s_mux_signals[3][0][22] ,
         \s_mux_signals[3][0][21] , \s_mux_signals[3][0][20] ,
         \s_mux_signals[3][0][19] , \s_mux_signals[3][0][18] ,
         \s_mux_signals[3][0][17] , \s_mux_signals[3][0][16] ,
         \s_mux_signals[3][0][15] , \s_mux_signals[3][0][14] ,
         \s_mux_signals[3][0][13] , \s_mux_signals[3][0][12] ,
         \s_mux_signals[3][0][11] , \s_mux_signals[3][0][10] ,
         \s_mux_signals[3][0][9] , \s_mux_signals[3][0][8] ,
         \s_mux_signals[3][0][7] , \s_mux_signals[3][0][6] ,
         \s_mux_signals[3][0][5] , \s_mux_signals[3][0][4] ,
         \s_mux_signals[3][0][3] , \s_mux_signals[3][0][2] ,
         \s_mux_signals[3][0][1] , \s_mux_signals[3][0][0] ,
         \s_mux_signals[3][8][31] , \s_mux_signals[3][8][30] ,
         \s_mux_signals[3][8][29] , \s_mux_signals[3][8][28] ,
         \s_mux_signals[3][8][27] , \s_mux_signals[3][8][26] ,
         \s_mux_signals[3][8][25] , \s_mux_signals[3][8][24] ,
         \s_mux_signals[3][8][23] , \s_mux_signals[3][8][22] ,
         \s_mux_signals[3][8][21] , \s_mux_signals[3][8][20] ,
         \s_mux_signals[3][8][19] , \s_mux_signals[3][8][18] ,
         \s_mux_signals[3][8][17] , \s_mux_signals[3][8][16] ,
         \s_mux_signals[3][8][15] , \s_mux_signals[3][8][14] ,
         \s_mux_signals[3][8][13] , \s_mux_signals[3][8][12] ,
         \s_mux_signals[3][8][11] , \s_mux_signals[3][8][10] ,
         \s_mux_signals[3][8][9] , \s_mux_signals[3][8][8] ,
         \s_mux_signals[3][8][7] , \s_mux_signals[3][8][6] ,
         \s_mux_signals[3][8][5] , \s_mux_signals[3][8][4] ,
         \s_mux_signals[3][8][3] , \s_mux_signals[3][8][2] ,
         \s_mux_signals[3][8][1] , \s_mux_signals[3][8][0] ,
         \s_mux_signals[3][16][31] , \s_mux_signals[3][16][30] ,
         \s_mux_signals[3][16][29] , \s_mux_signals[3][16][28] ,
         \s_mux_signals[3][16][27] , \s_mux_signals[3][16][26] ,
         \s_mux_signals[3][16][25] , \s_mux_signals[3][16][24] ,
         \s_mux_signals[3][16][23] , \s_mux_signals[3][16][22] ,
         \s_mux_signals[3][16][21] , \s_mux_signals[3][16][20] ,
         \s_mux_signals[3][16][19] , \s_mux_signals[3][16][18] ,
         \s_mux_signals[3][16][17] , \s_mux_signals[3][16][16] ,
         \s_mux_signals[3][16][15] , \s_mux_signals[3][16][14] ,
         \s_mux_signals[3][16][13] , \s_mux_signals[3][16][12] ,
         \s_mux_signals[3][16][11] , \s_mux_signals[3][16][10] ,
         \s_mux_signals[3][16][9] , \s_mux_signals[3][16][8] ,
         \s_mux_signals[3][16][7] , \s_mux_signals[3][16][6] ,
         \s_mux_signals[3][16][5] , \s_mux_signals[3][16][4] ,
         \s_mux_signals[3][16][3] , \s_mux_signals[3][16][2] ,
         \s_mux_signals[3][16][1] , \s_mux_signals[3][16][0] ,
         \s_mux_signals[3][24][31] , \s_mux_signals[3][24][30] ,
         \s_mux_signals[3][24][29] , \s_mux_signals[3][24][28] ,
         \s_mux_signals[3][24][27] , \s_mux_signals[3][24][26] ,
         \s_mux_signals[3][24][25] , \s_mux_signals[3][24][24] ,
         \s_mux_signals[3][24][23] , \s_mux_signals[3][24][22] ,
         \s_mux_signals[3][24][21] , \s_mux_signals[3][24][20] ,
         \s_mux_signals[3][24][19] , \s_mux_signals[3][24][18] ,
         \s_mux_signals[3][24][17] , \s_mux_signals[3][24][16] ,
         \s_mux_signals[3][24][15] , \s_mux_signals[3][24][14] ,
         \s_mux_signals[3][24][13] , \s_mux_signals[3][24][12] ,
         \s_mux_signals[3][24][11] , \s_mux_signals[3][24][10] ,
         \s_mux_signals[3][24][9] , \s_mux_signals[3][24][8] ,
         \s_mux_signals[3][24][7] , \s_mux_signals[3][24][6] ,
         \s_mux_signals[3][24][5] , \s_mux_signals[3][24][4] ,
         \s_mux_signals[3][24][3] , \s_mux_signals[3][24][2] ,
         \s_mux_signals[3][24][1] , \s_mux_signals[3][24][0] ,
         \s_mux_signals[4][0][31] , \s_mux_signals[4][0][30] ,
         \s_mux_signals[4][0][29] , \s_mux_signals[4][0][28] ,
         \s_mux_signals[4][0][27] , \s_mux_signals[4][0][26] ,
         \s_mux_signals[4][0][25] , \s_mux_signals[4][0][24] ,
         \s_mux_signals[4][0][23] , \s_mux_signals[4][0][22] ,
         \s_mux_signals[4][0][21] , \s_mux_signals[4][0][20] ,
         \s_mux_signals[4][0][19] , \s_mux_signals[4][0][18] ,
         \s_mux_signals[4][0][17] , \s_mux_signals[4][0][16] ,
         \s_mux_signals[4][0][15] , \s_mux_signals[4][0][14] ,
         \s_mux_signals[4][0][13] , \s_mux_signals[4][0][12] ,
         \s_mux_signals[4][0][11] , \s_mux_signals[4][0][10] ,
         \s_mux_signals[4][0][9] , \s_mux_signals[4][0][8] ,
         \s_mux_signals[4][0][7] , \s_mux_signals[4][0][6] ,
         \s_mux_signals[4][0][5] , \s_mux_signals[4][0][4] ,
         \s_mux_signals[4][0][3] , \s_mux_signals[4][0][2] ,
         \s_mux_signals[4][0][1] , \s_mux_signals[4][0][0] ,
         \s_mux_signals[4][16][31] , \s_mux_signals[4][16][30] ,
         \s_mux_signals[4][16][29] , \s_mux_signals[4][16][28] ,
         \s_mux_signals[4][16][27] , \s_mux_signals[4][16][26] ,
         \s_mux_signals[4][16][25] , \s_mux_signals[4][16][24] ,
         \s_mux_signals[4][16][23] , \s_mux_signals[4][16][22] ,
         \s_mux_signals[4][16][21] , \s_mux_signals[4][16][20] ,
         \s_mux_signals[4][16][19] , \s_mux_signals[4][16][18] ,
         \s_mux_signals[4][16][17] , \s_mux_signals[4][16][16] ,
         \s_mux_signals[4][16][15] , \s_mux_signals[4][16][14] ,
         \s_mux_signals[4][16][13] , \s_mux_signals[4][16][12] ,
         \s_mux_signals[4][16][11] , \s_mux_signals[4][16][10] ,
         \s_mux_signals[4][16][9] , \s_mux_signals[4][16][8] ,
         \s_mux_signals[4][16][7] , \s_mux_signals[4][16][6] ,
         \s_mux_signals[4][16][5] , \s_mux_signals[4][16][4] ,
         \s_mux_signals[4][16][3] , \s_mux_signals[4][16][2] ,
         \s_mux_signals[4][16][1] , \s_mux_signals[4][16][0] ,
         \s_mux_signals[5][0][31] , \s_mux_signals[5][0][30] ,
         \s_mux_signals[5][0][29] , \s_mux_signals[5][0][28] ,
         \s_mux_signals[5][0][27] , \s_mux_signals[5][0][26] ,
         \s_mux_signals[5][0][25] , \s_mux_signals[5][0][24] ,
         \s_mux_signals[5][0][23] , \s_mux_signals[5][0][22] ,
         \s_mux_signals[5][0][21] , \s_mux_signals[5][0][20] ,
         \s_mux_signals[5][0][19] , \s_mux_signals[5][0][18] ,
         \s_mux_signals[5][0][17] , \s_mux_signals[5][0][16] ,
         \s_mux_signals[5][0][15] , \s_mux_signals[5][0][14] ,
         \s_mux_signals[5][0][13] , \s_mux_signals[5][0][12] ,
         \s_mux_signals[5][0][11] , \s_mux_signals[5][0][10] ,
         \s_mux_signals[5][0][9] , \s_mux_signals[5][0][8] ,
         \s_mux_signals[5][0][7] , \s_mux_signals[5][0][6] ,
         \s_mux_signals[5][0][5] , \s_mux_signals[5][0][4] ,
         \s_mux_signals[5][0][3] , \s_mux_signals[5][0][2] ,
         \s_mux_signals[5][0][1] , \s_mux_signals[5][0][0] ,
         s_HIT_miss_Freg_Txor, s_sat_prediction_Toutput, s_btb_prediction, n1,
         n3, n5, n8, n6, n11, n12, n13, n14, n15, n16, n17, n18, n19, n20, n21,
         n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33, n34, n35,
         n36, n37, n38, n39, n40, n41, n42, n43, n44, n45, n46, n47, n48, n49,
         n50, n51, n52, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n224, n225,
         n226, n227, n228, n229, n230, n231, n232, n233, n234, n235, n236,
         n237, n238, n239, n240, n241, n242, n243, n244, n245, n246, n247,
         n248, n249, n250, n251, n252, n253, n254, n255, n256, n257, n258,
         n259, n260, n261, n262, n263, n264, n265, n266, n267, n268, n269,
         n270, n271, n272, n273, n274, n275, n276, n277, n278, n279, n280,
         n281, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n296, n297, n298, n299, n300, n301, n302,
         n303, n304, n305, n306, n307, n308, n309, n310, n311, n312, n313,
         n314, n315, n316, n317, n318, n319, n320, n321, n322, n323, n324,
         n325, n326, n327, n328, n329, n330, n331, n332, n333, n334, n335;
  wire   [31:0] s_cmpbits_Fcmp_Tencoder;
  wire   [4:0] s_selmuxes_Fencoder_Tmuxes;
  wire   [31:0] s_regenabl_entry;
  wire   [31:0] s_regenabl_target;
  wire   [31:0] s_regenabl_FrotateR_Tregs;
  wire   [31:0] s_regenabl_sat;
  wire   [31:0] s_updateSat_FregCmpBits_Tsats;
  wire   [31:0] s_prediction_Fsat_Tmuxes;
  assign n8 = BTB_enable;

  NComparatorWithEnable_NBIT32_0 NCmp_i_0 ( .A({n317, n314, n311, n308, n305, 
        n302, n299, n296, n293, n290, n287, n284, n281, n278, n275, n272, n269, 
        n266, n263, n260, n257, n254, n251, n248, n245, n242, n239, n236, n233, 
        n230, n227, n224}), .B({\s_entries_Freg_Tcmp[0][31] , 
        \s_entries_Freg_Tcmp[0][30] , \s_entries_Freg_Tcmp[0][29] , 
        \s_entries_Freg_Tcmp[0][28] , \s_entries_Freg_Tcmp[0][27] , 
        \s_entries_Freg_Tcmp[0][26] , \s_entries_Freg_Tcmp[0][25] , 
        \s_entries_Freg_Tcmp[0][24] , \s_entries_Freg_Tcmp[0][23] , 
        \s_entries_Freg_Tcmp[0][22] , \s_entries_Freg_Tcmp[0][21] , 
        \s_entries_Freg_Tcmp[0][20] , \s_entries_Freg_Tcmp[0][19] , 
        \s_entries_Freg_Tcmp[0][18] , \s_entries_Freg_Tcmp[0][17] , 
        \s_entries_Freg_Tcmp[0][16] , \s_entries_Freg_Tcmp[0][15] , 
        \s_entries_Freg_Tcmp[0][14] , \s_entries_Freg_Tcmp[0][13] , 
        \s_entries_Freg_Tcmp[0][12] , \s_entries_Freg_Tcmp[0][11] , 
        \s_entries_Freg_Tcmp[0][10] , \s_entries_Freg_Tcmp[0][9] , 
        \s_entries_Freg_Tcmp[0][8] , \s_entries_Freg_Tcmp[0][7] , 
        \s_entries_Freg_Tcmp[0][6] , \s_entries_Freg_Tcmp[0][5] , 
        \s_entries_Freg_Tcmp[0][4] , \s_entries_Freg_Tcmp[0][3] , 
        \s_entries_Freg_Tcmp[0][2] , \s_entries_Freg_Tcmp[0][1] , 
        \s_entries_Freg_Tcmp[0][0] }), .Enable(n321), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[0]) );
  NComparatorWithEnable_NBIT32_32 NCmp_i_1 ( .A({n315, n312, n309, n306, n303, 
        n300, n297, n294, n291, n288, n285, n282, n279, n276, n273, n270, n267, 
        n264, n261, n258, n255, n252, n249, n246, n243, n240, n237, n234, n231, 
        n228, n225, n222}), .B({\s_entries_Freg_Tcmp[1][31] , 
        \s_entries_Freg_Tcmp[1][30] , \s_entries_Freg_Tcmp[1][29] , 
        \s_entries_Freg_Tcmp[1][28] , \s_entries_Freg_Tcmp[1][27] , 
        \s_entries_Freg_Tcmp[1][26] , \s_entries_Freg_Tcmp[1][25] , 
        \s_entries_Freg_Tcmp[1][24] , \s_entries_Freg_Tcmp[1][23] , 
        \s_entries_Freg_Tcmp[1][22] , \s_entries_Freg_Tcmp[1][21] , 
        \s_entries_Freg_Tcmp[1][20] , \s_entries_Freg_Tcmp[1][19] , 
        \s_entries_Freg_Tcmp[1][18] , \s_entries_Freg_Tcmp[1][17] , 
        \s_entries_Freg_Tcmp[1][16] , \s_entries_Freg_Tcmp[1][15] , 
        \s_entries_Freg_Tcmp[1][14] , \s_entries_Freg_Tcmp[1][13] , 
        \s_entries_Freg_Tcmp[1][12] , \s_entries_Freg_Tcmp[1][11] , 
        \s_entries_Freg_Tcmp[1][10] , \s_entries_Freg_Tcmp[1][9] , 
        \s_entries_Freg_Tcmp[1][8] , \s_entries_Freg_Tcmp[1][7] , 
        \s_entries_Freg_Tcmp[1][6] , \s_entries_Freg_Tcmp[1][5] , 
        \s_entries_Freg_Tcmp[1][4] , \s_entries_Freg_Tcmp[1][3] , 
        \s_entries_Freg_Tcmp[1][2] , \s_entries_Freg_Tcmp[1][1] , 
        \s_entries_Freg_Tcmp[1][0] }), .Enable(n318), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[1]) );
  NComparatorWithEnable_NBIT32_31 NCmp_i_2 ( .A({n315, n312, n309, n306, n303, 
        n300, n297, n294, n291, n288, n285, n282, n279, n276, n273, n270, n267, 
        n264, n261, n258, n255, n252, n249, n246, n243, n240, n237, n234, n231, 
        n228, n225, n222}), .B({\s_entries_Freg_Tcmp[2][31] , 
        \s_entries_Freg_Tcmp[2][30] , \s_entries_Freg_Tcmp[2][29] , 
        \s_entries_Freg_Tcmp[2][28] , \s_entries_Freg_Tcmp[2][27] , 
        \s_entries_Freg_Tcmp[2][26] , \s_entries_Freg_Tcmp[2][25] , 
        \s_entries_Freg_Tcmp[2][24] , \s_entries_Freg_Tcmp[2][23] , 
        \s_entries_Freg_Tcmp[2][22] , \s_entries_Freg_Tcmp[2][21] , 
        \s_entries_Freg_Tcmp[2][20] , \s_entries_Freg_Tcmp[2][19] , 
        \s_entries_Freg_Tcmp[2][18] , \s_entries_Freg_Tcmp[2][17] , 
        \s_entries_Freg_Tcmp[2][16] , \s_entries_Freg_Tcmp[2][15] , 
        \s_entries_Freg_Tcmp[2][14] , \s_entries_Freg_Tcmp[2][13] , 
        \s_entries_Freg_Tcmp[2][12] , \s_entries_Freg_Tcmp[2][11] , 
        \s_entries_Freg_Tcmp[2][10] , \s_entries_Freg_Tcmp[2][9] , 
        \s_entries_Freg_Tcmp[2][8] , \s_entries_Freg_Tcmp[2][7] , 
        \s_entries_Freg_Tcmp[2][6] , \s_entries_Freg_Tcmp[2][5] , 
        \s_entries_Freg_Tcmp[2][4] , \s_entries_Freg_Tcmp[2][3] , 
        \s_entries_Freg_Tcmp[2][2] , \s_entries_Freg_Tcmp[2][1] , 
        \s_entries_Freg_Tcmp[2][0] }), .Enable(n323), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[2]) );
  NComparatorWithEnable_NBIT32_30 NCmp_i_3 ( .A({n315, n312, n309, n306, n303, 
        n300, n297, n294, n291, n288, n285, n282, n279, n276, n273, n270, n267, 
        n264, n261, n258, n255, n252, n249, n246, n243, n240, n237, n234, n231, 
        n228, n225, n222}), .B({\s_entries_Freg_Tcmp[3][31] , 
        \s_entries_Freg_Tcmp[3][30] , \s_entries_Freg_Tcmp[3][29] , 
        \s_entries_Freg_Tcmp[3][28] , \s_entries_Freg_Tcmp[3][27] , 
        \s_entries_Freg_Tcmp[3][26] , \s_entries_Freg_Tcmp[3][25] , 
        \s_entries_Freg_Tcmp[3][24] , \s_entries_Freg_Tcmp[3][23] , 
        \s_entries_Freg_Tcmp[3][22] , \s_entries_Freg_Tcmp[3][21] , 
        \s_entries_Freg_Tcmp[3][20] , \s_entries_Freg_Tcmp[3][19] , 
        \s_entries_Freg_Tcmp[3][18] , \s_entries_Freg_Tcmp[3][17] , 
        \s_entries_Freg_Tcmp[3][16] , \s_entries_Freg_Tcmp[3][15] , 
        \s_entries_Freg_Tcmp[3][14] , \s_entries_Freg_Tcmp[3][13] , 
        \s_entries_Freg_Tcmp[3][12] , \s_entries_Freg_Tcmp[3][11] , 
        \s_entries_Freg_Tcmp[3][10] , \s_entries_Freg_Tcmp[3][9] , 
        \s_entries_Freg_Tcmp[3][8] , \s_entries_Freg_Tcmp[3][7] , 
        \s_entries_Freg_Tcmp[3][6] , \s_entries_Freg_Tcmp[3][5] , 
        \s_entries_Freg_Tcmp[3][4] , \s_entries_Freg_Tcmp[3][3] , 
        \s_entries_Freg_Tcmp[3][2] , \s_entries_Freg_Tcmp[3][1] , 
        \s_entries_Freg_Tcmp[3][0] }), .Enable(n323), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[3]) );
  NComparatorWithEnable_NBIT32_29 NCmp_i_4 ( .A({n315, n312, n309, n306, n303, 
        n300, n297, n294, n291, n288, n285, n282, n279, n276, n273, n270, n267, 
        n264, n261, n258, n255, n252, n249, n246, n243, n240, n237, n234, n231, 
        n228, n225, n222}), .B({\s_entries_Freg_Tcmp[4][31] , 
        \s_entries_Freg_Tcmp[4][30] , \s_entries_Freg_Tcmp[4][29] , 
        \s_entries_Freg_Tcmp[4][28] , \s_entries_Freg_Tcmp[4][27] , 
        \s_entries_Freg_Tcmp[4][26] , \s_entries_Freg_Tcmp[4][25] , 
        \s_entries_Freg_Tcmp[4][24] , \s_entries_Freg_Tcmp[4][23] , 
        \s_entries_Freg_Tcmp[4][22] , \s_entries_Freg_Tcmp[4][21] , 
        \s_entries_Freg_Tcmp[4][20] , \s_entries_Freg_Tcmp[4][19] , 
        \s_entries_Freg_Tcmp[4][18] , \s_entries_Freg_Tcmp[4][17] , 
        \s_entries_Freg_Tcmp[4][16] , \s_entries_Freg_Tcmp[4][15] , 
        \s_entries_Freg_Tcmp[4][14] , \s_entries_Freg_Tcmp[4][13] , 
        \s_entries_Freg_Tcmp[4][12] , \s_entries_Freg_Tcmp[4][11] , 
        \s_entries_Freg_Tcmp[4][10] , \s_entries_Freg_Tcmp[4][9] , 
        \s_entries_Freg_Tcmp[4][8] , \s_entries_Freg_Tcmp[4][7] , 
        \s_entries_Freg_Tcmp[4][6] , \s_entries_Freg_Tcmp[4][5] , 
        \s_entries_Freg_Tcmp[4][4] , \s_entries_Freg_Tcmp[4][3] , 
        \s_entries_Freg_Tcmp[4][2] , \s_entries_Freg_Tcmp[4][1] , 
        \s_entries_Freg_Tcmp[4][0] }), .Enable(n323), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[4]) );
  NComparatorWithEnable_NBIT32_28 NCmp_i_5 ( .A({n315, n312, n309, n306, n303, 
        n300, n297, n294, n291, n288, n285, n282, n279, n276, n273, n270, n267, 
        n264, n261, n258, n255, n252, n249, n246, n243, n240, n237, n234, n231, 
        n228, n225, n222}), .B({\s_entries_Freg_Tcmp[5][31] , 
        \s_entries_Freg_Tcmp[5][30] , \s_entries_Freg_Tcmp[5][29] , 
        \s_entries_Freg_Tcmp[5][28] , \s_entries_Freg_Tcmp[5][27] , 
        \s_entries_Freg_Tcmp[5][26] , \s_entries_Freg_Tcmp[5][25] , 
        \s_entries_Freg_Tcmp[5][24] , \s_entries_Freg_Tcmp[5][23] , 
        \s_entries_Freg_Tcmp[5][22] , \s_entries_Freg_Tcmp[5][21] , 
        \s_entries_Freg_Tcmp[5][20] , \s_entries_Freg_Tcmp[5][19] , 
        \s_entries_Freg_Tcmp[5][18] , \s_entries_Freg_Tcmp[5][17] , 
        \s_entries_Freg_Tcmp[5][16] , \s_entries_Freg_Tcmp[5][15] , 
        \s_entries_Freg_Tcmp[5][14] , \s_entries_Freg_Tcmp[5][13] , 
        \s_entries_Freg_Tcmp[5][12] , \s_entries_Freg_Tcmp[5][11] , 
        \s_entries_Freg_Tcmp[5][10] , \s_entries_Freg_Tcmp[5][9] , 
        \s_entries_Freg_Tcmp[5][8] , \s_entries_Freg_Tcmp[5][7] , 
        \s_entries_Freg_Tcmp[5][6] , \s_entries_Freg_Tcmp[5][5] , 
        \s_entries_Freg_Tcmp[5][4] , \s_entries_Freg_Tcmp[5][3] , 
        \s_entries_Freg_Tcmp[5][2] , \s_entries_Freg_Tcmp[5][1] , 
        \s_entries_Freg_Tcmp[5][0] }), .Enable(n323), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[5]) );
  NComparatorWithEnable_NBIT32_27 NCmp_i_6 ( .A({n315, n312, n309, n306, n303, 
        n300, n297, n294, n291, n288, n285, n282, n279, n276, n273, n270, n267, 
        n264, n261, n258, n255, n252, n249, n246, n243, n240, n237, n234, n231, 
        n228, n225, n222}), .B({\s_entries_Freg_Tcmp[6][31] , 
        \s_entries_Freg_Tcmp[6][30] , \s_entries_Freg_Tcmp[6][29] , 
        \s_entries_Freg_Tcmp[6][28] , \s_entries_Freg_Tcmp[6][27] , 
        \s_entries_Freg_Tcmp[6][26] , \s_entries_Freg_Tcmp[6][25] , 
        \s_entries_Freg_Tcmp[6][24] , \s_entries_Freg_Tcmp[6][23] , 
        \s_entries_Freg_Tcmp[6][22] , \s_entries_Freg_Tcmp[6][21] , 
        \s_entries_Freg_Tcmp[6][20] , \s_entries_Freg_Tcmp[6][19] , 
        \s_entries_Freg_Tcmp[6][18] , \s_entries_Freg_Tcmp[6][17] , 
        \s_entries_Freg_Tcmp[6][16] , \s_entries_Freg_Tcmp[6][15] , 
        \s_entries_Freg_Tcmp[6][14] , \s_entries_Freg_Tcmp[6][13] , 
        \s_entries_Freg_Tcmp[6][12] , \s_entries_Freg_Tcmp[6][11] , 
        \s_entries_Freg_Tcmp[6][10] , \s_entries_Freg_Tcmp[6][9] , 
        \s_entries_Freg_Tcmp[6][8] , \s_entries_Freg_Tcmp[6][7] , 
        \s_entries_Freg_Tcmp[6][6] , \s_entries_Freg_Tcmp[6][5] , 
        \s_entries_Freg_Tcmp[6][4] , \s_entries_Freg_Tcmp[6][3] , 
        \s_entries_Freg_Tcmp[6][2] , \s_entries_Freg_Tcmp[6][1] , 
        \s_entries_Freg_Tcmp[6][0] }), .Enable(n323), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[6]) );
  NComparatorWithEnable_NBIT32_26 NCmp_i_7 ( .A({n315, n312, n309, n306, n303, 
        n300, n297, n294, n291, n288, n285, n282, n279, n276, n273, n270, n267, 
        n264, n261, n258, n255, n252, n249, n246, n243, n240, n237, n234, n231, 
        n228, n225, n222}), .B({\s_entries_Freg_Tcmp[7][31] , 
        \s_entries_Freg_Tcmp[7][30] , \s_entries_Freg_Tcmp[7][29] , 
        \s_entries_Freg_Tcmp[7][28] , \s_entries_Freg_Tcmp[7][27] , 
        \s_entries_Freg_Tcmp[7][26] , \s_entries_Freg_Tcmp[7][25] , 
        \s_entries_Freg_Tcmp[7][24] , \s_entries_Freg_Tcmp[7][23] , 
        \s_entries_Freg_Tcmp[7][22] , \s_entries_Freg_Tcmp[7][21] , 
        \s_entries_Freg_Tcmp[7][20] , \s_entries_Freg_Tcmp[7][19] , 
        \s_entries_Freg_Tcmp[7][18] , \s_entries_Freg_Tcmp[7][17] , 
        \s_entries_Freg_Tcmp[7][16] , \s_entries_Freg_Tcmp[7][15] , 
        \s_entries_Freg_Tcmp[7][14] , \s_entries_Freg_Tcmp[7][13] , 
        \s_entries_Freg_Tcmp[7][12] , \s_entries_Freg_Tcmp[7][11] , 
        \s_entries_Freg_Tcmp[7][10] , \s_entries_Freg_Tcmp[7][9] , 
        \s_entries_Freg_Tcmp[7][8] , \s_entries_Freg_Tcmp[7][7] , 
        \s_entries_Freg_Tcmp[7][6] , \s_entries_Freg_Tcmp[7][5] , 
        \s_entries_Freg_Tcmp[7][4] , \s_entries_Freg_Tcmp[7][3] , 
        \s_entries_Freg_Tcmp[7][2] , \s_entries_Freg_Tcmp[7][1] , 
        \s_entries_Freg_Tcmp[7][0] }), .Enable(n322), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[7]) );
  NComparatorWithEnable_NBIT32_25 NCmp_i_8 ( .A({n315, n312, n309, n306, n303, 
        n300, n297, n294, n291, n288, n285, n282, n279, n276, n273, n270, n267, 
        n264, n261, n258, n255, n252, n249, n246, n243, n240, n237, n234, n231, 
        n228, n225, n222}), .B({\s_entries_Freg_Tcmp[8][31] , 
        \s_entries_Freg_Tcmp[8][30] , \s_entries_Freg_Tcmp[8][29] , 
        \s_entries_Freg_Tcmp[8][28] , \s_entries_Freg_Tcmp[8][27] , 
        \s_entries_Freg_Tcmp[8][26] , \s_entries_Freg_Tcmp[8][25] , 
        \s_entries_Freg_Tcmp[8][24] , \s_entries_Freg_Tcmp[8][23] , 
        \s_entries_Freg_Tcmp[8][22] , \s_entries_Freg_Tcmp[8][21] , 
        \s_entries_Freg_Tcmp[8][20] , \s_entries_Freg_Tcmp[8][19] , 
        \s_entries_Freg_Tcmp[8][18] , \s_entries_Freg_Tcmp[8][17] , 
        \s_entries_Freg_Tcmp[8][16] , \s_entries_Freg_Tcmp[8][15] , 
        \s_entries_Freg_Tcmp[8][14] , \s_entries_Freg_Tcmp[8][13] , 
        \s_entries_Freg_Tcmp[8][12] , \s_entries_Freg_Tcmp[8][11] , 
        \s_entries_Freg_Tcmp[8][10] , \s_entries_Freg_Tcmp[8][9] , 
        \s_entries_Freg_Tcmp[8][8] , \s_entries_Freg_Tcmp[8][7] , 
        \s_entries_Freg_Tcmp[8][6] , \s_entries_Freg_Tcmp[8][5] , 
        \s_entries_Freg_Tcmp[8][4] , \s_entries_Freg_Tcmp[8][3] , 
        \s_entries_Freg_Tcmp[8][2] , \s_entries_Freg_Tcmp[8][1] , 
        \s_entries_Freg_Tcmp[8][0] }), .Enable(n322), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[8]) );
  NComparatorWithEnable_NBIT32_24 NCmp_i_9 ( .A({n315, n312, n309, n306, n303, 
        n300, n297, n294, n291, n288, n285, n282, n279, n276, n273, n270, n267, 
        n264, n261, n258, n255, n252, n249, n246, n243, n240, n237, n234, n231, 
        n228, n225, n222}), .B({\s_entries_Freg_Tcmp[9][31] , 
        \s_entries_Freg_Tcmp[9][30] , \s_entries_Freg_Tcmp[9][29] , 
        \s_entries_Freg_Tcmp[9][28] , \s_entries_Freg_Tcmp[9][27] , 
        \s_entries_Freg_Tcmp[9][26] , \s_entries_Freg_Tcmp[9][25] , 
        \s_entries_Freg_Tcmp[9][24] , \s_entries_Freg_Tcmp[9][23] , 
        \s_entries_Freg_Tcmp[9][22] , \s_entries_Freg_Tcmp[9][21] , 
        \s_entries_Freg_Tcmp[9][20] , \s_entries_Freg_Tcmp[9][19] , 
        \s_entries_Freg_Tcmp[9][18] , \s_entries_Freg_Tcmp[9][17] , 
        \s_entries_Freg_Tcmp[9][16] , \s_entries_Freg_Tcmp[9][15] , 
        \s_entries_Freg_Tcmp[9][14] , \s_entries_Freg_Tcmp[9][13] , 
        \s_entries_Freg_Tcmp[9][12] , \s_entries_Freg_Tcmp[9][11] , 
        \s_entries_Freg_Tcmp[9][10] , \s_entries_Freg_Tcmp[9][9] , 
        \s_entries_Freg_Tcmp[9][8] , \s_entries_Freg_Tcmp[9][7] , 
        \s_entries_Freg_Tcmp[9][6] , \s_entries_Freg_Tcmp[9][5] , 
        \s_entries_Freg_Tcmp[9][4] , \s_entries_Freg_Tcmp[9][3] , 
        \s_entries_Freg_Tcmp[9][2] , \s_entries_Freg_Tcmp[9][1] , 
        \s_entries_Freg_Tcmp[9][0] }), .Enable(n322), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[9]) );
  NComparatorWithEnable_NBIT32_23 NCmp_i_10 ( .A({n315, n312, n309, n306, n303, 
        n300, n297, n294, n291, n288, n285, n282, n279, n276, n273, n270, n267, 
        n264, n261, n258, n255, n252, n249, n246, n243, n240, n237, n234, n231, 
        n228, n225, n222}), .B({\s_entries_Freg_Tcmp[10][31] , 
        \s_entries_Freg_Tcmp[10][30] , \s_entries_Freg_Tcmp[10][29] , 
        \s_entries_Freg_Tcmp[10][28] , \s_entries_Freg_Tcmp[10][27] , 
        \s_entries_Freg_Tcmp[10][26] , \s_entries_Freg_Tcmp[10][25] , 
        \s_entries_Freg_Tcmp[10][24] , \s_entries_Freg_Tcmp[10][23] , 
        \s_entries_Freg_Tcmp[10][22] , \s_entries_Freg_Tcmp[10][21] , 
        \s_entries_Freg_Tcmp[10][20] , \s_entries_Freg_Tcmp[10][19] , 
        \s_entries_Freg_Tcmp[10][18] , \s_entries_Freg_Tcmp[10][17] , 
        \s_entries_Freg_Tcmp[10][16] , \s_entries_Freg_Tcmp[10][15] , 
        \s_entries_Freg_Tcmp[10][14] , \s_entries_Freg_Tcmp[10][13] , 
        \s_entries_Freg_Tcmp[10][12] , \s_entries_Freg_Tcmp[10][11] , 
        \s_entries_Freg_Tcmp[10][10] , \s_entries_Freg_Tcmp[10][9] , 
        \s_entries_Freg_Tcmp[10][8] , \s_entries_Freg_Tcmp[10][7] , 
        \s_entries_Freg_Tcmp[10][6] , \s_entries_Freg_Tcmp[10][5] , 
        \s_entries_Freg_Tcmp[10][4] , \s_entries_Freg_Tcmp[10][3] , 
        \s_entries_Freg_Tcmp[10][2] , \s_entries_Freg_Tcmp[10][1] , 
        \s_entries_Freg_Tcmp[10][0] }), .Enable(n322), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[10]) );
  NComparatorWithEnable_NBIT32_22 NCmp_i_11 ( .A({n315, n312, n309, n306, n303, 
        n300, n297, n294, n291, n288, n285, n282, n279, n276, n273, n270, n267, 
        n264, n261, n258, n255, n252, n249, n246, n243, n240, n237, n234, n231, 
        n228, n225, n222}), .B({\s_entries_Freg_Tcmp[11][31] , 
        \s_entries_Freg_Tcmp[11][30] , \s_entries_Freg_Tcmp[11][29] , 
        \s_entries_Freg_Tcmp[11][28] , \s_entries_Freg_Tcmp[11][27] , 
        \s_entries_Freg_Tcmp[11][26] , \s_entries_Freg_Tcmp[11][25] , 
        \s_entries_Freg_Tcmp[11][24] , \s_entries_Freg_Tcmp[11][23] , 
        \s_entries_Freg_Tcmp[11][22] , \s_entries_Freg_Tcmp[11][21] , 
        \s_entries_Freg_Tcmp[11][20] , \s_entries_Freg_Tcmp[11][19] , 
        \s_entries_Freg_Tcmp[11][18] , \s_entries_Freg_Tcmp[11][17] , 
        \s_entries_Freg_Tcmp[11][16] , \s_entries_Freg_Tcmp[11][15] , 
        \s_entries_Freg_Tcmp[11][14] , \s_entries_Freg_Tcmp[11][13] , 
        \s_entries_Freg_Tcmp[11][12] , \s_entries_Freg_Tcmp[11][11] , 
        \s_entries_Freg_Tcmp[11][10] , \s_entries_Freg_Tcmp[11][9] , 
        \s_entries_Freg_Tcmp[11][8] , \s_entries_Freg_Tcmp[11][7] , 
        \s_entries_Freg_Tcmp[11][6] , \s_entries_Freg_Tcmp[11][5] , 
        \s_entries_Freg_Tcmp[11][4] , \s_entries_Freg_Tcmp[11][3] , 
        \s_entries_Freg_Tcmp[11][2] , \s_entries_Freg_Tcmp[11][1] , 
        \s_entries_Freg_Tcmp[11][0] }), .Enable(n322), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[11]) );
  NComparatorWithEnable_NBIT32_21 NCmp_i_12 ( .A({n315, n312, n309, n306, n303, 
        n300, n297, n294, n291, n288, n285, n282, n279, n276, n273, n270, n267, 
        n264, n261, n258, n255, n252, n249, n246, n243, n240, n237, n234, n231, 
        n228, n225, n222}), .B({\s_entries_Freg_Tcmp[12][31] , 
        \s_entries_Freg_Tcmp[12][30] , \s_entries_Freg_Tcmp[12][29] , 
        \s_entries_Freg_Tcmp[12][28] , \s_entries_Freg_Tcmp[12][27] , 
        \s_entries_Freg_Tcmp[12][26] , \s_entries_Freg_Tcmp[12][25] , 
        \s_entries_Freg_Tcmp[12][24] , \s_entries_Freg_Tcmp[12][23] , 
        \s_entries_Freg_Tcmp[12][22] , \s_entries_Freg_Tcmp[12][21] , 
        \s_entries_Freg_Tcmp[12][20] , \s_entries_Freg_Tcmp[12][19] , 
        \s_entries_Freg_Tcmp[12][18] , \s_entries_Freg_Tcmp[12][17] , 
        \s_entries_Freg_Tcmp[12][16] , \s_entries_Freg_Tcmp[12][15] , 
        \s_entries_Freg_Tcmp[12][14] , \s_entries_Freg_Tcmp[12][13] , 
        \s_entries_Freg_Tcmp[12][12] , \s_entries_Freg_Tcmp[12][11] , 
        \s_entries_Freg_Tcmp[12][10] , \s_entries_Freg_Tcmp[12][9] , 
        \s_entries_Freg_Tcmp[12][8] , \s_entries_Freg_Tcmp[12][7] , 
        \s_entries_Freg_Tcmp[12][6] , \s_entries_Freg_Tcmp[12][5] , 
        \s_entries_Freg_Tcmp[12][4] , \s_entries_Freg_Tcmp[12][3] , 
        \s_entries_Freg_Tcmp[12][2] , \s_entries_Freg_Tcmp[12][1] , 
        \s_entries_Freg_Tcmp[12][0] }), .Enable(n322), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[12]) );
  NComparatorWithEnable_NBIT32_20 NCmp_i_13 ( .A({n316, n313, n310, n307, n304, 
        n301, n298, n295, n292, n289, n286, n283, n280, n277, n274, n271, n268, 
        n265, n262, n259, n256, n253, n250, n247, n244, n241, n238, n235, n232, 
        n229, n226, n223}), .B({\s_entries_Freg_Tcmp[13][31] , 
        \s_entries_Freg_Tcmp[13][30] , \s_entries_Freg_Tcmp[13][29] , 
        \s_entries_Freg_Tcmp[13][28] , \s_entries_Freg_Tcmp[13][27] , 
        \s_entries_Freg_Tcmp[13][26] , \s_entries_Freg_Tcmp[13][25] , 
        \s_entries_Freg_Tcmp[13][24] , \s_entries_Freg_Tcmp[13][23] , 
        \s_entries_Freg_Tcmp[13][22] , \s_entries_Freg_Tcmp[13][21] , 
        \s_entries_Freg_Tcmp[13][20] , \s_entries_Freg_Tcmp[13][19] , 
        \s_entries_Freg_Tcmp[13][18] , \s_entries_Freg_Tcmp[13][17] , 
        \s_entries_Freg_Tcmp[13][16] , \s_entries_Freg_Tcmp[13][15] , 
        \s_entries_Freg_Tcmp[13][14] , \s_entries_Freg_Tcmp[13][13] , 
        \s_entries_Freg_Tcmp[13][12] , \s_entries_Freg_Tcmp[13][11] , 
        \s_entries_Freg_Tcmp[13][10] , \s_entries_Freg_Tcmp[13][9] , 
        \s_entries_Freg_Tcmp[13][8] , \s_entries_Freg_Tcmp[13][7] , 
        \s_entries_Freg_Tcmp[13][6] , \s_entries_Freg_Tcmp[13][5] , 
        \s_entries_Freg_Tcmp[13][4] , \s_entries_Freg_Tcmp[13][3] , 
        \s_entries_Freg_Tcmp[13][2] , \s_entries_Freg_Tcmp[13][1] , 
        \s_entries_Freg_Tcmp[13][0] }), .Enable(n321), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[13]) );
  NComparatorWithEnable_NBIT32_19 NCmp_i_14 ( .A({n316, n313, n310, n307, n304, 
        n301, n298, n295, n292, n289, n286, n283, n280, n277, n274, n271, n268, 
        n265, n262, n259, n256, n253, n250, n247, n244, n241, n238, n235, n232, 
        n229, n226, n223}), .B({\s_entries_Freg_Tcmp[14][31] , 
        \s_entries_Freg_Tcmp[14][30] , \s_entries_Freg_Tcmp[14][29] , 
        \s_entries_Freg_Tcmp[14][28] , \s_entries_Freg_Tcmp[14][27] , 
        \s_entries_Freg_Tcmp[14][26] , \s_entries_Freg_Tcmp[14][25] , 
        \s_entries_Freg_Tcmp[14][24] , \s_entries_Freg_Tcmp[14][23] , 
        \s_entries_Freg_Tcmp[14][22] , \s_entries_Freg_Tcmp[14][21] , 
        \s_entries_Freg_Tcmp[14][20] , \s_entries_Freg_Tcmp[14][19] , 
        \s_entries_Freg_Tcmp[14][18] , \s_entries_Freg_Tcmp[14][17] , 
        \s_entries_Freg_Tcmp[14][16] , \s_entries_Freg_Tcmp[14][15] , 
        \s_entries_Freg_Tcmp[14][14] , \s_entries_Freg_Tcmp[14][13] , 
        \s_entries_Freg_Tcmp[14][12] , \s_entries_Freg_Tcmp[14][11] , 
        \s_entries_Freg_Tcmp[14][10] , \s_entries_Freg_Tcmp[14][9] , 
        \s_entries_Freg_Tcmp[14][8] , \s_entries_Freg_Tcmp[14][7] , 
        \s_entries_Freg_Tcmp[14][6] , \s_entries_Freg_Tcmp[14][5] , 
        \s_entries_Freg_Tcmp[14][4] , \s_entries_Freg_Tcmp[14][3] , 
        \s_entries_Freg_Tcmp[14][2] , \s_entries_Freg_Tcmp[14][1] , 
        \s_entries_Freg_Tcmp[14][0] }), .Enable(n321), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[14]) );
  NComparatorWithEnable_NBIT32_18 NCmp_i_15 ( .A({n316, n313, n310, n307, n304, 
        n301, n298, n295, n292, n289, n286, n283, n280, n277, n274, n271, n268, 
        n265, n262, n259, n256, n253, n250, n247, n244, n241, n238, n235, n232, 
        n229, n226, n223}), .B({\s_entries_Freg_Tcmp[15][31] , 
        \s_entries_Freg_Tcmp[15][30] , \s_entries_Freg_Tcmp[15][29] , 
        \s_entries_Freg_Tcmp[15][28] , \s_entries_Freg_Tcmp[15][27] , 
        \s_entries_Freg_Tcmp[15][26] , \s_entries_Freg_Tcmp[15][25] , 
        \s_entries_Freg_Tcmp[15][24] , \s_entries_Freg_Tcmp[15][23] , 
        \s_entries_Freg_Tcmp[15][22] , \s_entries_Freg_Tcmp[15][21] , 
        \s_entries_Freg_Tcmp[15][20] , \s_entries_Freg_Tcmp[15][19] , 
        \s_entries_Freg_Tcmp[15][18] , \s_entries_Freg_Tcmp[15][17] , 
        \s_entries_Freg_Tcmp[15][16] , \s_entries_Freg_Tcmp[15][15] , 
        \s_entries_Freg_Tcmp[15][14] , \s_entries_Freg_Tcmp[15][13] , 
        \s_entries_Freg_Tcmp[15][12] , \s_entries_Freg_Tcmp[15][11] , 
        \s_entries_Freg_Tcmp[15][10] , \s_entries_Freg_Tcmp[15][9] , 
        \s_entries_Freg_Tcmp[15][8] , \s_entries_Freg_Tcmp[15][7] , 
        \s_entries_Freg_Tcmp[15][6] , \s_entries_Freg_Tcmp[15][5] , 
        \s_entries_Freg_Tcmp[15][4] , \s_entries_Freg_Tcmp[15][3] , 
        \s_entries_Freg_Tcmp[15][2] , \s_entries_Freg_Tcmp[15][1] , 
        \s_entries_Freg_Tcmp[15][0] }), .Enable(n321), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[15]) );
  NComparatorWithEnable_NBIT32_17 NCmp_i_16 ( .A({n316, n313, n310, n307, n304, 
        n301, n298, n295, n292, n289, n286, n283, n280, n277, n274, n271, n268, 
        n265, n262, n259, n256, n253, n250, n247, n244, n241, n238, n235, n232, 
        n229, n226, n223}), .B({\s_entries_Freg_Tcmp[16][31] , 
        \s_entries_Freg_Tcmp[16][30] , \s_entries_Freg_Tcmp[16][29] , 
        \s_entries_Freg_Tcmp[16][28] , \s_entries_Freg_Tcmp[16][27] , 
        \s_entries_Freg_Tcmp[16][26] , \s_entries_Freg_Tcmp[16][25] , 
        \s_entries_Freg_Tcmp[16][24] , \s_entries_Freg_Tcmp[16][23] , 
        \s_entries_Freg_Tcmp[16][22] , \s_entries_Freg_Tcmp[16][21] , 
        \s_entries_Freg_Tcmp[16][20] , \s_entries_Freg_Tcmp[16][19] , 
        \s_entries_Freg_Tcmp[16][18] , \s_entries_Freg_Tcmp[16][17] , 
        \s_entries_Freg_Tcmp[16][16] , \s_entries_Freg_Tcmp[16][15] , 
        \s_entries_Freg_Tcmp[16][14] , \s_entries_Freg_Tcmp[16][13] , 
        \s_entries_Freg_Tcmp[16][12] , \s_entries_Freg_Tcmp[16][11] , 
        \s_entries_Freg_Tcmp[16][10] , \s_entries_Freg_Tcmp[16][9] , 
        \s_entries_Freg_Tcmp[16][8] , \s_entries_Freg_Tcmp[16][7] , 
        \s_entries_Freg_Tcmp[16][6] , \s_entries_Freg_Tcmp[16][5] , 
        \s_entries_Freg_Tcmp[16][4] , \s_entries_Freg_Tcmp[16][3] , 
        \s_entries_Freg_Tcmp[16][2] , \s_entries_Freg_Tcmp[16][1] , 
        \s_entries_Freg_Tcmp[16][0] }), .Enable(n321), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[16]) );
  NComparatorWithEnable_NBIT32_16 NCmp_i_17 ( .A({n316, n313, n310, n307, n304, 
        n301, n298, n295, n292, n289, n286, n283, n280, n277, n274, n271, n268, 
        n265, n262, n259, n256, n253, n250, n247, n244, n241, n238, n235, n232, 
        n229, n226, n223}), .B({\s_entries_Freg_Tcmp[17][31] , 
        \s_entries_Freg_Tcmp[17][30] , \s_entries_Freg_Tcmp[17][29] , 
        \s_entries_Freg_Tcmp[17][28] , \s_entries_Freg_Tcmp[17][27] , 
        \s_entries_Freg_Tcmp[17][26] , \s_entries_Freg_Tcmp[17][25] , 
        \s_entries_Freg_Tcmp[17][24] , \s_entries_Freg_Tcmp[17][23] , 
        \s_entries_Freg_Tcmp[17][22] , \s_entries_Freg_Tcmp[17][21] , 
        \s_entries_Freg_Tcmp[17][20] , \s_entries_Freg_Tcmp[17][19] , 
        \s_entries_Freg_Tcmp[17][18] , \s_entries_Freg_Tcmp[17][17] , 
        \s_entries_Freg_Tcmp[17][16] , \s_entries_Freg_Tcmp[17][15] , 
        \s_entries_Freg_Tcmp[17][14] , \s_entries_Freg_Tcmp[17][13] , 
        \s_entries_Freg_Tcmp[17][12] , \s_entries_Freg_Tcmp[17][11] , 
        \s_entries_Freg_Tcmp[17][10] , \s_entries_Freg_Tcmp[17][9] , 
        \s_entries_Freg_Tcmp[17][8] , \s_entries_Freg_Tcmp[17][7] , 
        \s_entries_Freg_Tcmp[17][6] , \s_entries_Freg_Tcmp[17][5] , 
        \s_entries_Freg_Tcmp[17][4] , \s_entries_Freg_Tcmp[17][3] , 
        \s_entries_Freg_Tcmp[17][2] , \s_entries_Freg_Tcmp[17][1] , 
        \s_entries_Freg_Tcmp[17][0] }), .Enable(n321), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[17]) );
  NComparatorWithEnable_NBIT32_15 NCmp_i_18 ( .A({n316, n313, n310, n307, n304, 
        n301, n298, n295, n292, n289, n286, n283, n280, n277, n274, n271, n268, 
        n265, n262, n259, n256, n253, n250, n247, n244, n241, n238, n235, n232, 
        n229, n226, n223}), .B({\s_entries_Freg_Tcmp[18][31] , 
        \s_entries_Freg_Tcmp[18][30] , \s_entries_Freg_Tcmp[18][29] , 
        \s_entries_Freg_Tcmp[18][28] , \s_entries_Freg_Tcmp[18][27] , 
        \s_entries_Freg_Tcmp[18][26] , \s_entries_Freg_Tcmp[18][25] , 
        \s_entries_Freg_Tcmp[18][24] , \s_entries_Freg_Tcmp[18][23] , 
        \s_entries_Freg_Tcmp[18][22] , \s_entries_Freg_Tcmp[18][21] , 
        \s_entries_Freg_Tcmp[18][20] , \s_entries_Freg_Tcmp[18][19] , 
        \s_entries_Freg_Tcmp[18][18] , \s_entries_Freg_Tcmp[18][17] , 
        \s_entries_Freg_Tcmp[18][16] , \s_entries_Freg_Tcmp[18][15] , 
        \s_entries_Freg_Tcmp[18][14] , \s_entries_Freg_Tcmp[18][13] , 
        \s_entries_Freg_Tcmp[18][12] , \s_entries_Freg_Tcmp[18][11] , 
        \s_entries_Freg_Tcmp[18][10] , \s_entries_Freg_Tcmp[18][9] , 
        \s_entries_Freg_Tcmp[18][8] , \s_entries_Freg_Tcmp[18][7] , 
        \s_entries_Freg_Tcmp[18][6] , \s_entries_Freg_Tcmp[18][5] , 
        \s_entries_Freg_Tcmp[18][4] , \s_entries_Freg_Tcmp[18][3] , 
        \s_entries_Freg_Tcmp[18][2] , \s_entries_Freg_Tcmp[18][1] , 
        \s_entries_Freg_Tcmp[18][0] }), .Enable(n320), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[18]) );
  NComparatorWithEnable_NBIT32_14 NCmp_i_19 ( .A({n316, n313, n310, n307, n304, 
        n301, n298, n295, n292, n289, n286, n283, n280, n277, n274, n271, n268, 
        n265, n262, n259, n256, n253, n250, n247, n244, n241, n238, n235, n232, 
        n229, n226, n223}), .B({\s_entries_Freg_Tcmp[19][31] , 
        \s_entries_Freg_Tcmp[19][30] , \s_entries_Freg_Tcmp[19][29] , 
        \s_entries_Freg_Tcmp[19][28] , \s_entries_Freg_Tcmp[19][27] , 
        \s_entries_Freg_Tcmp[19][26] , \s_entries_Freg_Tcmp[19][25] , 
        \s_entries_Freg_Tcmp[19][24] , \s_entries_Freg_Tcmp[19][23] , 
        \s_entries_Freg_Tcmp[19][22] , \s_entries_Freg_Tcmp[19][21] , 
        \s_entries_Freg_Tcmp[19][20] , \s_entries_Freg_Tcmp[19][19] , 
        \s_entries_Freg_Tcmp[19][18] , \s_entries_Freg_Tcmp[19][17] , 
        \s_entries_Freg_Tcmp[19][16] , \s_entries_Freg_Tcmp[19][15] , 
        \s_entries_Freg_Tcmp[19][14] , \s_entries_Freg_Tcmp[19][13] , 
        \s_entries_Freg_Tcmp[19][12] , \s_entries_Freg_Tcmp[19][11] , 
        \s_entries_Freg_Tcmp[19][10] , \s_entries_Freg_Tcmp[19][9] , 
        \s_entries_Freg_Tcmp[19][8] , \s_entries_Freg_Tcmp[19][7] , 
        \s_entries_Freg_Tcmp[19][6] , \s_entries_Freg_Tcmp[19][5] , 
        \s_entries_Freg_Tcmp[19][4] , \s_entries_Freg_Tcmp[19][3] , 
        \s_entries_Freg_Tcmp[19][2] , \s_entries_Freg_Tcmp[19][1] , 
        \s_entries_Freg_Tcmp[19][0] }), .Enable(n320), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[19]) );
  NComparatorWithEnable_NBIT32_13 NCmp_i_20 ( .A({n316, n313, n310, n307, n304, 
        n301, n298, n295, n292, n289, n286, n283, n280, n277, n274, n271, n268, 
        n265, n262, n259, n256, n253, n250, n247, n244, n241, n238, n235, n232, 
        n229, n226, n223}), .B({\s_entries_Freg_Tcmp[20][31] , 
        \s_entries_Freg_Tcmp[20][30] , \s_entries_Freg_Tcmp[20][29] , 
        \s_entries_Freg_Tcmp[20][28] , \s_entries_Freg_Tcmp[20][27] , 
        \s_entries_Freg_Tcmp[20][26] , \s_entries_Freg_Tcmp[20][25] , 
        \s_entries_Freg_Tcmp[20][24] , \s_entries_Freg_Tcmp[20][23] , 
        \s_entries_Freg_Tcmp[20][22] , \s_entries_Freg_Tcmp[20][21] , 
        \s_entries_Freg_Tcmp[20][20] , \s_entries_Freg_Tcmp[20][19] , 
        \s_entries_Freg_Tcmp[20][18] , \s_entries_Freg_Tcmp[20][17] , 
        \s_entries_Freg_Tcmp[20][16] , \s_entries_Freg_Tcmp[20][15] , 
        \s_entries_Freg_Tcmp[20][14] , \s_entries_Freg_Tcmp[20][13] , 
        \s_entries_Freg_Tcmp[20][12] , \s_entries_Freg_Tcmp[20][11] , 
        \s_entries_Freg_Tcmp[20][10] , \s_entries_Freg_Tcmp[20][9] , 
        \s_entries_Freg_Tcmp[20][8] , \s_entries_Freg_Tcmp[20][7] , 
        \s_entries_Freg_Tcmp[20][6] , \s_entries_Freg_Tcmp[20][5] , 
        \s_entries_Freg_Tcmp[20][4] , \s_entries_Freg_Tcmp[20][3] , 
        \s_entries_Freg_Tcmp[20][2] , \s_entries_Freg_Tcmp[20][1] , 
        \s_entries_Freg_Tcmp[20][0] }), .Enable(n320), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[20]) );
  NComparatorWithEnable_NBIT32_12 NCmp_i_21 ( .A({n316, n313, n310, n307, n304, 
        n301, n298, n295, n292, n289, n286, n283, n280, n277, n274, n271, n268, 
        n265, n262, n259, n256, n253, n250, n247, n244, n241, n238, n235, n232, 
        n229, n226, n223}), .B({\s_entries_Freg_Tcmp[21][31] , 
        \s_entries_Freg_Tcmp[21][30] , \s_entries_Freg_Tcmp[21][29] , 
        \s_entries_Freg_Tcmp[21][28] , \s_entries_Freg_Tcmp[21][27] , 
        \s_entries_Freg_Tcmp[21][26] , \s_entries_Freg_Tcmp[21][25] , 
        \s_entries_Freg_Tcmp[21][24] , \s_entries_Freg_Tcmp[21][23] , 
        \s_entries_Freg_Tcmp[21][22] , \s_entries_Freg_Tcmp[21][21] , 
        \s_entries_Freg_Tcmp[21][20] , \s_entries_Freg_Tcmp[21][19] , 
        \s_entries_Freg_Tcmp[21][18] , \s_entries_Freg_Tcmp[21][17] , 
        \s_entries_Freg_Tcmp[21][16] , \s_entries_Freg_Tcmp[21][15] , 
        \s_entries_Freg_Tcmp[21][14] , \s_entries_Freg_Tcmp[21][13] , 
        \s_entries_Freg_Tcmp[21][12] , \s_entries_Freg_Tcmp[21][11] , 
        \s_entries_Freg_Tcmp[21][10] , \s_entries_Freg_Tcmp[21][9] , 
        \s_entries_Freg_Tcmp[21][8] , \s_entries_Freg_Tcmp[21][7] , 
        \s_entries_Freg_Tcmp[21][6] , \s_entries_Freg_Tcmp[21][5] , 
        \s_entries_Freg_Tcmp[21][4] , \s_entries_Freg_Tcmp[21][3] , 
        \s_entries_Freg_Tcmp[21][2] , \s_entries_Freg_Tcmp[21][1] , 
        \s_entries_Freg_Tcmp[21][0] }), .Enable(n320), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[21]) );
  NComparatorWithEnable_NBIT32_11 NCmp_i_22 ( .A({n316, n313, n310, n307, n304, 
        n301, n298, n295, n292, n289, n286, n283, n280, n277, n274, n271, n268, 
        n265, n262, n259, n256, n253, n250, n247, n244, n241, n238, n235, n232, 
        n229, n226, n223}), .B({\s_entries_Freg_Tcmp[22][31] , 
        \s_entries_Freg_Tcmp[22][30] , \s_entries_Freg_Tcmp[22][29] , 
        \s_entries_Freg_Tcmp[22][28] , \s_entries_Freg_Tcmp[22][27] , 
        \s_entries_Freg_Tcmp[22][26] , \s_entries_Freg_Tcmp[22][25] , 
        \s_entries_Freg_Tcmp[22][24] , \s_entries_Freg_Tcmp[22][23] , 
        \s_entries_Freg_Tcmp[22][22] , \s_entries_Freg_Tcmp[22][21] , 
        \s_entries_Freg_Tcmp[22][20] , \s_entries_Freg_Tcmp[22][19] , 
        \s_entries_Freg_Tcmp[22][18] , \s_entries_Freg_Tcmp[22][17] , 
        \s_entries_Freg_Tcmp[22][16] , \s_entries_Freg_Tcmp[22][15] , 
        \s_entries_Freg_Tcmp[22][14] , \s_entries_Freg_Tcmp[22][13] , 
        \s_entries_Freg_Tcmp[22][12] , \s_entries_Freg_Tcmp[22][11] , 
        \s_entries_Freg_Tcmp[22][10] , \s_entries_Freg_Tcmp[22][9] , 
        \s_entries_Freg_Tcmp[22][8] , \s_entries_Freg_Tcmp[22][7] , 
        \s_entries_Freg_Tcmp[22][6] , \s_entries_Freg_Tcmp[22][5] , 
        \s_entries_Freg_Tcmp[22][4] , \s_entries_Freg_Tcmp[22][3] , 
        \s_entries_Freg_Tcmp[22][2] , \s_entries_Freg_Tcmp[22][1] , 
        \s_entries_Freg_Tcmp[22][0] }), .Enable(n320), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[22]) );
  NComparatorWithEnable_NBIT32_10 NCmp_i_23 ( .A({n316, n313, n310, n307, n304, 
        n301, n298, n295, n292, n289, n286, n283, n280, n277, n274, n271, n268, 
        n265, n262, n259, n256, n253, n250, n247, n244, n241, n238, n235, n232, 
        n229, n226, n223}), .B({\s_entries_Freg_Tcmp[23][31] , 
        \s_entries_Freg_Tcmp[23][30] , \s_entries_Freg_Tcmp[23][29] , 
        \s_entries_Freg_Tcmp[23][28] , \s_entries_Freg_Tcmp[23][27] , 
        \s_entries_Freg_Tcmp[23][26] , \s_entries_Freg_Tcmp[23][25] , 
        \s_entries_Freg_Tcmp[23][24] , \s_entries_Freg_Tcmp[23][23] , 
        \s_entries_Freg_Tcmp[23][22] , \s_entries_Freg_Tcmp[23][21] , 
        \s_entries_Freg_Tcmp[23][20] , \s_entries_Freg_Tcmp[23][19] , 
        \s_entries_Freg_Tcmp[23][18] , \s_entries_Freg_Tcmp[23][17] , 
        \s_entries_Freg_Tcmp[23][16] , \s_entries_Freg_Tcmp[23][15] , 
        \s_entries_Freg_Tcmp[23][14] , \s_entries_Freg_Tcmp[23][13] , 
        \s_entries_Freg_Tcmp[23][12] , \s_entries_Freg_Tcmp[23][11] , 
        \s_entries_Freg_Tcmp[23][10] , \s_entries_Freg_Tcmp[23][9] , 
        \s_entries_Freg_Tcmp[23][8] , \s_entries_Freg_Tcmp[23][7] , 
        \s_entries_Freg_Tcmp[23][6] , \s_entries_Freg_Tcmp[23][5] , 
        \s_entries_Freg_Tcmp[23][4] , \s_entries_Freg_Tcmp[23][3] , 
        \s_entries_Freg_Tcmp[23][2] , \s_entries_Freg_Tcmp[23][1] , 
        \s_entries_Freg_Tcmp[23][0] }), .Enable(n320), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[23]) );
  NComparatorWithEnable_NBIT32_9 NCmp_i_24 ( .A({n316, n313, n310, n307, n304, 
        n301, n298, n295, n292, n289, n286, n283, n280, n277, n274, n271, n268, 
        n265, n262, n259, n256, n253, n250, n247, n244, n241, n238, n235, n232, 
        n229, n226, n223}), .B({\s_entries_Freg_Tcmp[24][31] , 
        \s_entries_Freg_Tcmp[24][30] , \s_entries_Freg_Tcmp[24][29] , 
        \s_entries_Freg_Tcmp[24][28] , \s_entries_Freg_Tcmp[24][27] , 
        \s_entries_Freg_Tcmp[24][26] , \s_entries_Freg_Tcmp[24][25] , 
        \s_entries_Freg_Tcmp[24][24] , \s_entries_Freg_Tcmp[24][23] , 
        \s_entries_Freg_Tcmp[24][22] , \s_entries_Freg_Tcmp[24][21] , 
        \s_entries_Freg_Tcmp[24][20] , \s_entries_Freg_Tcmp[24][19] , 
        \s_entries_Freg_Tcmp[24][18] , \s_entries_Freg_Tcmp[24][17] , 
        \s_entries_Freg_Tcmp[24][16] , \s_entries_Freg_Tcmp[24][15] , 
        \s_entries_Freg_Tcmp[24][14] , \s_entries_Freg_Tcmp[24][13] , 
        \s_entries_Freg_Tcmp[24][12] , \s_entries_Freg_Tcmp[24][11] , 
        \s_entries_Freg_Tcmp[24][10] , \s_entries_Freg_Tcmp[24][9] , 
        \s_entries_Freg_Tcmp[24][8] , \s_entries_Freg_Tcmp[24][7] , 
        \s_entries_Freg_Tcmp[24][6] , \s_entries_Freg_Tcmp[24][5] , 
        \s_entries_Freg_Tcmp[24][4] , \s_entries_Freg_Tcmp[24][3] , 
        \s_entries_Freg_Tcmp[24][2] , \s_entries_Freg_Tcmp[24][1] , 
        \s_entries_Freg_Tcmp[24][0] }), .Enable(n319), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[24]) );
  NComparatorWithEnable_NBIT32_8 NCmp_i_25 ( .A({n317, n314, n311, n308, n305, 
        n302, n299, n296, n293, n290, n287, n284, n281, n278, n275, n272, n269, 
        n266, n263, n260, n257, n254, n251, n248, n245, n242, n239, n236, n233, 
        n230, n227, n224}), .B({\s_entries_Freg_Tcmp[25][31] , 
        \s_entries_Freg_Tcmp[25][30] , \s_entries_Freg_Tcmp[25][29] , 
        \s_entries_Freg_Tcmp[25][28] , \s_entries_Freg_Tcmp[25][27] , 
        \s_entries_Freg_Tcmp[25][26] , \s_entries_Freg_Tcmp[25][25] , 
        \s_entries_Freg_Tcmp[25][24] , \s_entries_Freg_Tcmp[25][23] , 
        \s_entries_Freg_Tcmp[25][22] , \s_entries_Freg_Tcmp[25][21] , 
        \s_entries_Freg_Tcmp[25][20] , \s_entries_Freg_Tcmp[25][19] , 
        \s_entries_Freg_Tcmp[25][18] , \s_entries_Freg_Tcmp[25][17] , 
        \s_entries_Freg_Tcmp[25][16] , \s_entries_Freg_Tcmp[25][15] , 
        \s_entries_Freg_Tcmp[25][14] , \s_entries_Freg_Tcmp[25][13] , 
        \s_entries_Freg_Tcmp[25][12] , \s_entries_Freg_Tcmp[25][11] , 
        \s_entries_Freg_Tcmp[25][10] , \s_entries_Freg_Tcmp[25][9] , 
        \s_entries_Freg_Tcmp[25][8] , \s_entries_Freg_Tcmp[25][7] , 
        \s_entries_Freg_Tcmp[25][6] , \s_entries_Freg_Tcmp[25][5] , 
        \s_entries_Freg_Tcmp[25][4] , \s_entries_Freg_Tcmp[25][3] , 
        \s_entries_Freg_Tcmp[25][2] , \s_entries_Freg_Tcmp[25][1] , 
        \s_entries_Freg_Tcmp[25][0] }), .Enable(n319), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[25]) );
  NComparatorWithEnable_NBIT32_7 NCmp_i_26 ( .A({n317, n314, n311, n308, n305, 
        n302, n299, n296, n293, n290, n287, n284, n281, n278, n275, n272, n269, 
        n266, n263, n260, n257, n254, n251, n248, n245, n242, n239, n236, n233, 
        n230, n227, n224}), .B({\s_entries_Freg_Tcmp[26][31] , 
        \s_entries_Freg_Tcmp[26][30] , \s_entries_Freg_Tcmp[26][29] , 
        \s_entries_Freg_Tcmp[26][28] , \s_entries_Freg_Tcmp[26][27] , 
        \s_entries_Freg_Tcmp[26][26] , \s_entries_Freg_Tcmp[26][25] , 
        \s_entries_Freg_Tcmp[26][24] , \s_entries_Freg_Tcmp[26][23] , 
        \s_entries_Freg_Tcmp[26][22] , \s_entries_Freg_Tcmp[26][21] , 
        \s_entries_Freg_Tcmp[26][20] , \s_entries_Freg_Tcmp[26][19] , 
        \s_entries_Freg_Tcmp[26][18] , \s_entries_Freg_Tcmp[26][17] , 
        \s_entries_Freg_Tcmp[26][16] , \s_entries_Freg_Tcmp[26][15] , 
        \s_entries_Freg_Tcmp[26][14] , \s_entries_Freg_Tcmp[26][13] , 
        \s_entries_Freg_Tcmp[26][12] , \s_entries_Freg_Tcmp[26][11] , 
        \s_entries_Freg_Tcmp[26][10] , \s_entries_Freg_Tcmp[26][9] , 
        \s_entries_Freg_Tcmp[26][8] , \s_entries_Freg_Tcmp[26][7] , 
        \s_entries_Freg_Tcmp[26][6] , \s_entries_Freg_Tcmp[26][5] , 
        \s_entries_Freg_Tcmp[26][4] , \s_entries_Freg_Tcmp[26][3] , 
        \s_entries_Freg_Tcmp[26][2] , \s_entries_Freg_Tcmp[26][1] , 
        \s_entries_Freg_Tcmp[26][0] }), .Enable(n319), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[26]) );
  NComparatorWithEnable_NBIT32_6 NCmp_i_27 ( .A({n317, n314, n311, n308, n305, 
        n302, n299, n296, n293, n290, n287, n284, n281, n278, n275, n272, n269, 
        n266, n263, n260, n257, n254, n251, n248, n245, n242, n239, n236, n233, 
        n230, n227, n224}), .B({\s_entries_Freg_Tcmp[27][31] , 
        \s_entries_Freg_Tcmp[27][30] , \s_entries_Freg_Tcmp[27][29] , 
        \s_entries_Freg_Tcmp[27][28] , \s_entries_Freg_Tcmp[27][27] , 
        \s_entries_Freg_Tcmp[27][26] , \s_entries_Freg_Tcmp[27][25] , 
        \s_entries_Freg_Tcmp[27][24] , \s_entries_Freg_Tcmp[27][23] , 
        \s_entries_Freg_Tcmp[27][22] , \s_entries_Freg_Tcmp[27][21] , 
        \s_entries_Freg_Tcmp[27][20] , \s_entries_Freg_Tcmp[27][19] , 
        \s_entries_Freg_Tcmp[27][18] , \s_entries_Freg_Tcmp[27][17] , 
        \s_entries_Freg_Tcmp[27][16] , \s_entries_Freg_Tcmp[27][15] , 
        \s_entries_Freg_Tcmp[27][14] , \s_entries_Freg_Tcmp[27][13] , 
        \s_entries_Freg_Tcmp[27][12] , \s_entries_Freg_Tcmp[27][11] , 
        \s_entries_Freg_Tcmp[27][10] , \s_entries_Freg_Tcmp[27][9] , 
        \s_entries_Freg_Tcmp[27][8] , \s_entries_Freg_Tcmp[27][7] , 
        \s_entries_Freg_Tcmp[27][6] , \s_entries_Freg_Tcmp[27][5] , 
        \s_entries_Freg_Tcmp[27][4] , \s_entries_Freg_Tcmp[27][3] , 
        \s_entries_Freg_Tcmp[27][2] , \s_entries_Freg_Tcmp[27][1] , 
        \s_entries_Freg_Tcmp[27][0] }), .Enable(n319), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[27]) );
  NComparatorWithEnable_NBIT32_5 NCmp_i_28 ( .A({n317, n314, n311, n308, n305, 
        n302, n299, n296, n293, n290, n287, n284, n281, n278, n275, n272, n269, 
        n266, n263, n260, n257, n254, n251, n248, n245, n242, n239, n236, n233, 
        n230, n227, n224}), .B({\s_entries_Freg_Tcmp[28][31] , 
        \s_entries_Freg_Tcmp[28][30] , \s_entries_Freg_Tcmp[28][29] , 
        \s_entries_Freg_Tcmp[28][28] , \s_entries_Freg_Tcmp[28][27] , 
        \s_entries_Freg_Tcmp[28][26] , \s_entries_Freg_Tcmp[28][25] , 
        \s_entries_Freg_Tcmp[28][24] , \s_entries_Freg_Tcmp[28][23] , 
        \s_entries_Freg_Tcmp[28][22] , \s_entries_Freg_Tcmp[28][21] , 
        \s_entries_Freg_Tcmp[28][20] , \s_entries_Freg_Tcmp[28][19] , 
        \s_entries_Freg_Tcmp[28][18] , \s_entries_Freg_Tcmp[28][17] , 
        \s_entries_Freg_Tcmp[28][16] , \s_entries_Freg_Tcmp[28][15] , 
        \s_entries_Freg_Tcmp[28][14] , \s_entries_Freg_Tcmp[28][13] , 
        \s_entries_Freg_Tcmp[28][12] , \s_entries_Freg_Tcmp[28][11] , 
        \s_entries_Freg_Tcmp[28][10] , \s_entries_Freg_Tcmp[28][9] , 
        \s_entries_Freg_Tcmp[28][8] , \s_entries_Freg_Tcmp[28][7] , 
        \s_entries_Freg_Tcmp[28][6] , \s_entries_Freg_Tcmp[28][5] , 
        \s_entries_Freg_Tcmp[28][4] , \s_entries_Freg_Tcmp[28][3] , 
        \s_entries_Freg_Tcmp[28][2] , \s_entries_Freg_Tcmp[28][1] , 
        \s_entries_Freg_Tcmp[28][0] }), .Enable(n319), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[28]) );
  NComparatorWithEnable_NBIT32_4 NCmp_i_29 ( .A({n317, n314, n311, n308, n305, 
        n302, n299, n296, n293, n290, n287, n284, n281, n278, n275, n272, n269, 
        n266, n263, n260, n257, n254, n251, n248, n245, n242, n239, n236, n233, 
        n230, n227, n224}), .B({\s_entries_Freg_Tcmp[29][31] , 
        \s_entries_Freg_Tcmp[29][30] , \s_entries_Freg_Tcmp[29][29] , 
        \s_entries_Freg_Tcmp[29][28] , \s_entries_Freg_Tcmp[29][27] , 
        \s_entries_Freg_Tcmp[29][26] , \s_entries_Freg_Tcmp[29][25] , 
        \s_entries_Freg_Tcmp[29][24] , \s_entries_Freg_Tcmp[29][23] , 
        \s_entries_Freg_Tcmp[29][22] , \s_entries_Freg_Tcmp[29][21] , 
        \s_entries_Freg_Tcmp[29][20] , \s_entries_Freg_Tcmp[29][19] , 
        \s_entries_Freg_Tcmp[29][18] , \s_entries_Freg_Tcmp[29][17] , 
        \s_entries_Freg_Tcmp[29][16] , \s_entries_Freg_Tcmp[29][15] , 
        \s_entries_Freg_Tcmp[29][14] , \s_entries_Freg_Tcmp[29][13] , 
        \s_entries_Freg_Tcmp[29][12] , \s_entries_Freg_Tcmp[29][11] , 
        \s_entries_Freg_Tcmp[29][10] , \s_entries_Freg_Tcmp[29][9] , 
        \s_entries_Freg_Tcmp[29][8] , \s_entries_Freg_Tcmp[29][7] , 
        \s_entries_Freg_Tcmp[29][6] , \s_entries_Freg_Tcmp[29][5] , 
        \s_entries_Freg_Tcmp[29][4] , \s_entries_Freg_Tcmp[29][3] , 
        \s_entries_Freg_Tcmp[29][2] , \s_entries_Freg_Tcmp[29][1] , 
        \s_entries_Freg_Tcmp[29][0] }), .Enable(n319), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[29]) );
  NComparatorWithEnable_NBIT32_3 NCmp_i_30 ( .A({n317, n314, n311, n308, n305, 
        n302, n299, n296, n293, n290, n287, n284, n281, n278, n275, n272, n269, 
        n266, n263, n260, n257, n254, n251, n248, n245, n242, n239, n236, n233, 
        n230, n227, n224}), .B({\s_entries_Freg_Tcmp[30][31] , 
        \s_entries_Freg_Tcmp[30][30] , \s_entries_Freg_Tcmp[30][29] , 
        \s_entries_Freg_Tcmp[30][28] , \s_entries_Freg_Tcmp[30][27] , 
        \s_entries_Freg_Tcmp[30][26] , \s_entries_Freg_Tcmp[30][25] , 
        \s_entries_Freg_Tcmp[30][24] , \s_entries_Freg_Tcmp[30][23] , 
        \s_entries_Freg_Tcmp[30][22] , \s_entries_Freg_Tcmp[30][21] , 
        \s_entries_Freg_Tcmp[30][20] , \s_entries_Freg_Tcmp[30][19] , 
        \s_entries_Freg_Tcmp[30][18] , \s_entries_Freg_Tcmp[30][17] , 
        \s_entries_Freg_Tcmp[30][16] , \s_entries_Freg_Tcmp[30][15] , 
        \s_entries_Freg_Tcmp[30][14] , \s_entries_Freg_Tcmp[30][13] , 
        \s_entries_Freg_Tcmp[30][12] , \s_entries_Freg_Tcmp[30][11] , 
        \s_entries_Freg_Tcmp[30][10] , \s_entries_Freg_Tcmp[30][9] , 
        \s_entries_Freg_Tcmp[30][8] , \s_entries_Freg_Tcmp[30][7] , 
        \s_entries_Freg_Tcmp[30][6] , \s_entries_Freg_Tcmp[30][5] , 
        \s_entries_Freg_Tcmp[30][4] , \s_entries_Freg_Tcmp[30][3] , 
        \s_entries_Freg_Tcmp[30][2] , \s_entries_Freg_Tcmp[30][1] , 
        \s_entries_Freg_Tcmp[30][0] }), .Enable(n318), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[30]) );
  NComparatorWithEnable_NBIT32_2 NCmp_i_31 ( .A({n317, n314, n311, n308, n305, 
        n302, n299, n296, n293, n290, n287, n284, n281, n278, n275, n272, n269, 
        n266, n263, n260, n257, n254, n251, n248, n245, n242, n239, n236, n233, 
        n230, n227, n224}), .B({\s_entries_Freg_Tcmp[31][31] , 
        \s_entries_Freg_Tcmp[31][30] , \s_entries_Freg_Tcmp[31][29] , 
        \s_entries_Freg_Tcmp[31][28] , \s_entries_Freg_Tcmp[31][27] , 
        \s_entries_Freg_Tcmp[31][26] , \s_entries_Freg_Tcmp[31][25] , 
        \s_entries_Freg_Tcmp[31][24] , \s_entries_Freg_Tcmp[31][23] , 
        \s_entries_Freg_Tcmp[31][22] , \s_entries_Freg_Tcmp[31][21] , 
        \s_entries_Freg_Tcmp[31][20] , \s_entries_Freg_Tcmp[31][19] , 
        \s_entries_Freg_Tcmp[31][18] , \s_entries_Freg_Tcmp[31][17] , 
        \s_entries_Freg_Tcmp[31][16] , \s_entries_Freg_Tcmp[31][15] , 
        \s_entries_Freg_Tcmp[31][14] , \s_entries_Freg_Tcmp[31][13] , 
        \s_entries_Freg_Tcmp[31][12] , \s_entries_Freg_Tcmp[31][11] , 
        \s_entries_Freg_Tcmp[31][10] , \s_entries_Freg_Tcmp[31][9] , 
        \s_entries_Freg_Tcmp[31][8] , \s_entries_Freg_Tcmp[31][7] , 
        \s_entries_Freg_Tcmp[31][6] , \s_entries_Freg_Tcmp[31][5] , 
        \s_entries_Freg_Tcmp[31][4] , \s_entries_Freg_Tcmp[31][3] , 
        \s_entries_Freg_Tcmp[31][2] , \s_entries_Freg_Tcmp[31][1] , 
        \s_entries_Freg_Tcmp[31][0] }), .Enable(n318), .ComparatorBit(
        s_cmpbits_Fcmp_Tencoder[31]) );
  ORGate_NX1_N32_0 ORGate32X1 ( .A(s_cmpbits_Fcmp_Tencoder), .B({1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .Y(s_HIT_miss) );
  NPriorityEncoder_NBIT_OUT5 PriorityEncoder32X5 ( .data_in(
        s_cmpbits_Fcmp_Tencoder), .enable(n322), .data_out({
        s_selmuxes_Fencoder_Tmuxes[4:1], n5}) );
  NRegister_N32_107 EntrReg_i_0 ( .clk(BTB_clk), .reset(n333), .data_in({n219, 
        n216, n213, n210, n207, n204, n201, n198, n195, n192, n189, n186, n183, 
        n180, n177, n174, n171, n168, n165, n162, n159, n156, n153, n150, n147, 
        n144, n141, n138, n135, n132, n129, n126}), .enable(n17), .load(
        s_regenabl_entry[31]), .data_out({\s_entries_Freg_Tcmp[0][31] , 
        \s_entries_Freg_Tcmp[0][30] , \s_entries_Freg_Tcmp[0][29] , 
        \s_entries_Freg_Tcmp[0][28] , \s_entries_Freg_Tcmp[0][27] , 
        \s_entries_Freg_Tcmp[0][26] , \s_entries_Freg_Tcmp[0][25] , 
        \s_entries_Freg_Tcmp[0][24] , \s_entries_Freg_Tcmp[0][23] , 
        \s_entries_Freg_Tcmp[0][22] , \s_entries_Freg_Tcmp[0][21] , 
        \s_entries_Freg_Tcmp[0][20] , \s_entries_Freg_Tcmp[0][19] , 
        \s_entries_Freg_Tcmp[0][18] , \s_entries_Freg_Tcmp[0][17] , 
        \s_entries_Freg_Tcmp[0][16] , \s_entries_Freg_Tcmp[0][15] , 
        \s_entries_Freg_Tcmp[0][14] , \s_entries_Freg_Tcmp[0][13] , 
        \s_entries_Freg_Tcmp[0][12] , \s_entries_Freg_Tcmp[0][11] , 
        \s_entries_Freg_Tcmp[0][10] , \s_entries_Freg_Tcmp[0][9] , 
        \s_entries_Freg_Tcmp[0][8] , \s_entries_Freg_Tcmp[0][7] , 
        \s_entries_Freg_Tcmp[0][6] , \s_entries_Freg_Tcmp[0][5] , 
        \s_entries_Freg_Tcmp[0][4] , \s_entries_Freg_Tcmp[0][3] , 
        \s_entries_Freg_Tcmp[0][2] , \s_entries_Freg_Tcmp[0][1] , 
        \s_entries_Freg_Tcmp[0][0] }) );
  NRegister_N32_106 EntrReg_i_1 ( .clk(BTB_clk), .reset(n333), .data_in({n219, 
        n216, n213, n210, n207, n204, n201, n198, n195, n192, n189, n186, n183, 
        n180, n177, n174, n171, n168, n165, n162, n159, n156, n153, n150, n147, 
        n144, n141, n138, n135, n132, n129, n126}), .enable(n17), .load(
        s_regenabl_entry[30]), .data_out({\s_entries_Freg_Tcmp[1][31] , 
        \s_entries_Freg_Tcmp[1][30] , \s_entries_Freg_Tcmp[1][29] , 
        \s_entries_Freg_Tcmp[1][28] , \s_entries_Freg_Tcmp[1][27] , 
        \s_entries_Freg_Tcmp[1][26] , \s_entries_Freg_Tcmp[1][25] , 
        \s_entries_Freg_Tcmp[1][24] , \s_entries_Freg_Tcmp[1][23] , 
        \s_entries_Freg_Tcmp[1][22] , \s_entries_Freg_Tcmp[1][21] , 
        \s_entries_Freg_Tcmp[1][20] , \s_entries_Freg_Tcmp[1][19] , 
        \s_entries_Freg_Tcmp[1][18] , \s_entries_Freg_Tcmp[1][17] , 
        \s_entries_Freg_Tcmp[1][16] , \s_entries_Freg_Tcmp[1][15] , 
        \s_entries_Freg_Tcmp[1][14] , \s_entries_Freg_Tcmp[1][13] , 
        \s_entries_Freg_Tcmp[1][12] , \s_entries_Freg_Tcmp[1][11] , 
        \s_entries_Freg_Tcmp[1][10] , \s_entries_Freg_Tcmp[1][9] , 
        \s_entries_Freg_Tcmp[1][8] , \s_entries_Freg_Tcmp[1][7] , 
        \s_entries_Freg_Tcmp[1][6] , \s_entries_Freg_Tcmp[1][5] , 
        \s_entries_Freg_Tcmp[1][4] , \s_entries_Freg_Tcmp[1][3] , 
        \s_entries_Freg_Tcmp[1][2] , \s_entries_Freg_Tcmp[1][1] , 
        \s_entries_Freg_Tcmp[1][0] }) );
  NRegister_N32_105 EntrReg_i_2 ( .clk(BTB_clk), .reset(n332), .data_in({n219, 
        n216, n213, n210, n207, n204, n201, n198, n195, n192, n189, n186, n183, 
        n180, n177, n174, n171, n168, n165, n162, n159, n156, n153, n150, n147, 
        n144, n141, n138, n135, n132, n129, n126}), .enable(n17), .load(
        s_regenabl_entry[29]), .data_out({\s_entries_Freg_Tcmp[2][31] , 
        \s_entries_Freg_Tcmp[2][30] , \s_entries_Freg_Tcmp[2][29] , 
        \s_entries_Freg_Tcmp[2][28] , \s_entries_Freg_Tcmp[2][27] , 
        \s_entries_Freg_Tcmp[2][26] , \s_entries_Freg_Tcmp[2][25] , 
        \s_entries_Freg_Tcmp[2][24] , \s_entries_Freg_Tcmp[2][23] , 
        \s_entries_Freg_Tcmp[2][22] , \s_entries_Freg_Tcmp[2][21] , 
        \s_entries_Freg_Tcmp[2][20] , \s_entries_Freg_Tcmp[2][19] , 
        \s_entries_Freg_Tcmp[2][18] , \s_entries_Freg_Tcmp[2][17] , 
        \s_entries_Freg_Tcmp[2][16] , \s_entries_Freg_Tcmp[2][15] , 
        \s_entries_Freg_Tcmp[2][14] , \s_entries_Freg_Tcmp[2][13] , 
        \s_entries_Freg_Tcmp[2][12] , \s_entries_Freg_Tcmp[2][11] , 
        \s_entries_Freg_Tcmp[2][10] , \s_entries_Freg_Tcmp[2][9] , 
        \s_entries_Freg_Tcmp[2][8] , \s_entries_Freg_Tcmp[2][7] , 
        \s_entries_Freg_Tcmp[2][6] , \s_entries_Freg_Tcmp[2][5] , 
        \s_entries_Freg_Tcmp[2][4] , \s_entries_Freg_Tcmp[2][3] , 
        \s_entries_Freg_Tcmp[2][2] , \s_entries_Freg_Tcmp[2][1] , 
        \s_entries_Freg_Tcmp[2][0] }) );
  NRegister_N32_104 EntrReg_i_3 ( .clk(BTB_clk), .reset(n333), .data_in({n219, 
        n216, n213, n210, n207, n204, n201, n198, n195, n192, n189, n186, n183, 
        n180, n177, n174, n171, n168, n165, n162, n159, n156, n153, n150, n147, 
        n144, n141, n138, n135, n132, n129, n126}), .enable(n17), .load(
        s_regenabl_entry[28]), .data_out({\s_entries_Freg_Tcmp[3][31] , 
        \s_entries_Freg_Tcmp[3][30] , \s_entries_Freg_Tcmp[3][29] , 
        \s_entries_Freg_Tcmp[3][28] , \s_entries_Freg_Tcmp[3][27] , 
        \s_entries_Freg_Tcmp[3][26] , \s_entries_Freg_Tcmp[3][25] , 
        \s_entries_Freg_Tcmp[3][24] , \s_entries_Freg_Tcmp[3][23] , 
        \s_entries_Freg_Tcmp[3][22] , \s_entries_Freg_Tcmp[3][21] , 
        \s_entries_Freg_Tcmp[3][20] , \s_entries_Freg_Tcmp[3][19] , 
        \s_entries_Freg_Tcmp[3][18] , \s_entries_Freg_Tcmp[3][17] , 
        \s_entries_Freg_Tcmp[3][16] , \s_entries_Freg_Tcmp[3][15] , 
        \s_entries_Freg_Tcmp[3][14] , \s_entries_Freg_Tcmp[3][13] , 
        \s_entries_Freg_Tcmp[3][12] , \s_entries_Freg_Tcmp[3][11] , 
        \s_entries_Freg_Tcmp[3][10] , \s_entries_Freg_Tcmp[3][9] , 
        \s_entries_Freg_Tcmp[3][8] , \s_entries_Freg_Tcmp[3][7] , 
        \s_entries_Freg_Tcmp[3][6] , \s_entries_Freg_Tcmp[3][5] , 
        \s_entries_Freg_Tcmp[3][4] , \s_entries_Freg_Tcmp[3][3] , 
        \s_entries_Freg_Tcmp[3][2] , \s_entries_Freg_Tcmp[3][1] , 
        \s_entries_Freg_Tcmp[3][0] }) );
  NRegister_N32_103 EntrReg_i_4 ( .clk(BTB_clk), .reset(n333), .data_in({n219, 
        n216, n213, n210, n207, n204, n201, n198, n195, n192, n189, n186, n183, 
        n180, n177, n174, n171, n168, n165, n162, n159, n156, n153, n150, n147, 
        n144, n141, n138, n135, n132, n129, n126}), .enable(n17), .load(
        s_regenabl_entry[27]), .data_out({\s_entries_Freg_Tcmp[4][31] , 
        \s_entries_Freg_Tcmp[4][30] , \s_entries_Freg_Tcmp[4][29] , 
        \s_entries_Freg_Tcmp[4][28] , \s_entries_Freg_Tcmp[4][27] , 
        \s_entries_Freg_Tcmp[4][26] , \s_entries_Freg_Tcmp[4][25] , 
        \s_entries_Freg_Tcmp[4][24] , \s_entries_Freg_Tcmp[4][23] , 
        \s_entries_Freg_Tcmp[4][22] , \s_entries_Freg_Tcmp[4][21] , 
        \s_entries_Freg_Tcmp[4][20] , \s_entries_Freg_Tcmp[4][19] , 
        \s_entries_Freg_Tcmp[4][18] , \s_entries_Freg_Tcmp[4][17] , 
        \s_entries_Freg_Tcmp[4][16] , \s_entries_Freg_Tcmp[4][15] , 
        \s_entries_Freg_Tcmp[4][14] , \s_entries_Freg_Tcmp[4][13] , 
        \s_entries_Freg_Tcmp[4][12] , \s_entries_Freg_Tcmp[4][11] , 
        \s_entries_Freg_Tcmp[4][10] , \s_entries_Freg_Tcmp[4][9] , 
        \s_entries_Freg_Tcmp[4][8] , \s_entries_Freg_Tcmp[4][7] , 
        \s_entries_Freg_Tcmp[4][6] , \s_entries_Freg_Tcmp[4][5] , 
        \s_entries_Freg_Tcmp[4][4] , \s_entries_Freg_Tcmp[4][3] , 
        \s_entries_Freg_Tcmp[4][2] , \s_entries_Freg_Tcmp[4][1] , 
        \s_entries_Freg_Tcmp[4][0] }) );
  NRegister_N32_102 EntrReg_i_5 ( .clk(BTB_clk), .reset(n333), .data_in({n219, 
        n216, n213, n210, n207, n204, n201, n198, n195, n192, n189, n186, n183, 
        n180, n177, n174, n171, n168, n165, n162, n159, n156, n153, n150, n147, 
        n144, n141, n138, n135, n132, n129, n126}), .enable(n17), .load(
        s_regenabl_entry[26]), .data_out({\s_entries_Freg_Tcmp[5][31] , 
        \s_entries_Freg_Tcmp[5][30] , \s_entries_Freg_Tcmp[5][29] , 
        \s_entries_Freg_Tcmp[5][28] , \s_entries_Freg_Tcmp[5][27] , 
        \s_entries_Freg_Tcmp[5][26] , \s_entries_Freg_Tcmp[5][25] , 
        \s_entries_Freg_Tcmp[5][24] , \s_entries_Freg_Tcmp[5][23] , 
        \s_entries_Freg_Tcmp[5][22] , \s_entries_Freg_Tcmp[5][21] , 
        \s_entries_Freg_Tcmp[5][20] , \s_entries_Freg_Tcmp[5][19] , 
        \s_entries_Freg_Tcmp[5][18] , \s_entries_Freg_Tcmp[5][17] , 
        \s_entries_Freg_Tcmp[5][16] , \s_entries_Freg_Tcmp[5][15] , 
        \s_entries_Freg_Tcmp[5][14] , \s_entries_Freg_Tcmp[5][13] , 
        \s_entries_Freg_Tcmp[5][12] , \s_entries_Freg_Tcmp[5][11] , 
        \s_entries_Freg_Tcmp[5][10] , \s_entries_Freg_Tcmp[5][9] , 
        \s_entries_Freg_Tcmp[5][8] , \s_entries_Freg_Tcmp[5][7] , 
        \s_entries_Freg_Tcmp[5][6] , \s_entries_Freg_Tcmp[5][5] , 
        \s_entries_Freg_Tcmp[5][4] , \s_entries_Freg_Tcmp[5][3] , 
        \s_entries_Freg_Tcmp[5][2] , \s_entries_Freg_Tcmp[5][1] , 
        \s_entries_Freg_Tcmp[5][0] }) );
  NRegister_N32_101 EntrReg_i_6 ( .clk(BTB_clk), .reset(n332), .data_in({n219, 
        n216, n213, n210, n207, n204, n201, n198, n195, n192, n189, n186, n183, 
        n180, n177, n174, n171, n168, n165, n162, n159, n156, n153, n150, n147, 
        n144, n141, n138, n135, n132, n129, n126}), .enable(n17), .load(
        s_regenabl_entry[25]), .data_out({\s_entries_Freg_Tcmp[6][31] , 
        \s_entries_Freg_Tcmp[6][30] , \s_entries_Freg_Tcmp[6][29] , 
        \s_entries_Freg_Tcmp[6][28] , \s_entries_Freg_Tcmp[6][27] , 
        \s_entries_Freg_Tcmp[6][26] , \s_entries_Freg_Tcmp[6][25] , 
        \s_entries_Freg_Tcmp[6][24] , \s_entries_Freg_Tcmp[6][23] , 
        \s_entries_Freg_Tcmp[6][22] , \s_entries_Freg_Tcmp[6][21] , 
        \s_entries_Freg_Tcmp[6][20] , \s_entries_Freg_Tcmp[6][19] , 
        \s_entries_Freg_Tcmp[6][18] , \s_entries_Freg_Tcmp[6][17] , 
        \s_entries_Freg_Tcmp[6][16] , \s_entries_Freg_Tcmp[6][15] , 
        \s_entries_Freg_Tcmp[6][14] , \s_entries_Freg_Tcmp[6][13] , 
        \s_entries_Freg_Tcmp[6][12] , \s_entries_Freg_Tcmp[6][11] , 
        \s_entries_Freg_Tcmp[6][10] , \s_entries_Freg_Tcmp[6][9] , 
        \s_entries_Freg_Tcmp[6][8] , \s_entries_Freg_Tcmp[6][7] , 
        \s_entries_Freg_Tcmp[6][6] , \s_entries_Freg_Tcmp[6][5] , 
        \s_entries_Freg_Tcmp[6][4] , \s_entries_Freg_Tcmp[6][3] , 
        \s_entries_Freg_Tcmp[6][2] , \s_entries_Freg_Tcmp[6][1] , 
        \s_entries_Freg_Tcmp[6][0] }) );
  NRegister_N32_100 EntrReg_i_7 ( .clk(BTB_clk), .reset(n332), .data_in({n219, 
        n216, n213, n210, n207, n204, n201, n198, n195, n192, n189, n186, n183, 
        n180, n177, n174, n171, n168, n165, n162, n159, n156, n153, n150, n147, 
        n144, n141, n138, n135, n132, n129, n126}), .enable(n17), .load(
        s_regenabl_entry[24]), .data_out({\s_entries_Freg_Tcmp[7][31] , 
        \s_entries_Freg_Tcmp[7][30] , \s_entries_Freg_Tcmp[7][29] , 
        \s_entries_Freg_Tcmp[7][28] , \s_entries_Freg_Tcmp[7][27] , 
        \s_entries_Freg_Tcmp[7][26] , \s_entries_Freg_Tcmp[7][25] , 
        \s_entries_Freg_Tcmp[7][24] , \s_entries_Freg_Tcmp[7][23] , 
        \s_entries_Freg_Tcmp[7][22] , \s_entries_Freg_Tcmp[7][21] , 
        \s_entries_Freg_Tcmp[7][20] , \s_entries_Freg_Tcmp[7][19] , 
        \s_entries_Freg_Tcmp[7][18] , \s_entries_Freg_Tcmp[7][17] , 
        \s_entries_Freg_Tcmp[7][16] , \s_entries_Freg_Tcmp[7][15] , 
        \s_entries_Freg_Tcmp[7][14] , \s_entries_Freg_Tcmp[7][13] , 
        \s_entries_Freg_Tcmp[7][12] , \s_entries_Freg_Tcmp[7][11] , 
        \s_entries_Freg_Tcmp[7][10] , \s_entries_Freg_Tcmp[7][9] , 
        \s_entries_Freg_Tcmp[7][8] , \s_entries_Freg_Tcmp[7][7] , 
        \s_entries_Freg_Tcmp[7][6] , \s_entries_Freg_Tcmp[7][5] , 
        \s_entries_Freg_Tcmp[7][4] , \s_entries_Freg_Tcmp[7][3] , 
        \s_entries_Freg_Tcmp[7][2] , \s_entries_Freg_Tcmp[7][1] , 
        \s_entries_Freg_Tcmp[7][0] }) );
  NRegister_N32_99 EntrReg_i_8 ( .clk(BTB_clk), .reset(n332), .data_in({n219, 
        n216, n213, n210, n207, n204, n201, n198, n195, n192, n189, n186, n183, 
        n180, n177, n174, n171, n168, n165, n162, n159, n156, n153, n150, n147, 
        n144, n141, n138, n135, n132, n129, n126}), .enable(n17), .load(
        s_regenabl_entry[23]), .data_out({\s_entries_Freg_Tcmp[8][31] , 
        \s_entries_Freg_Tcmp[8][30] , \s_entries_Freg_Tcmp[8][29] , 
        \s_entries_Freg_Tcmp[8][28] , \s_entries_Freg_Tcmp[8][27] , 
        \s_entries_Freg_Tcmp[8][26] , \s_entries_Freg_Tcmp[8][25] , 
        \s_entries_Freg_Tcmp[8][24] , \s_entries_Freg_Tcmp[8][23] , 
        \s_entries_Freg_Tcmp[8][22] , \s_entries_Freg_Tcmp[8][21] , 
        \s_entries_Freg_Tcmp[8][20] , \s_entries_Freg_Tcmp[8][19] , 
        \s_entries_Freg_Tcmp[8][18] , \s_entries_Freg_Tcmp[8][17] , 
        \s_entries_Freg_Tcmp[8][16] , \s_entries_Freg_Tcmp[8][15] , 
        \s_entries_Freg_Tcmp[8][14] , \s_entries_Freg_Tcmp[8][13] , 
        \s_entries_Freg_Tcmp[8][12] , \s_entries_Freg_Tcmp[8][11] , 
        \s_entries_Freg_Tcmp[8][10] , \s_entries_Freg_Tcmp[8][9] , 
        \s_entries_Freg_Tcmp[8][8] , \s_entries_Freg_Tcmp[8][7] , 
        \s_entries_Freg_Tcmp[8][6] , \s_entries_Freg_Tcmp[8][5] , 
        \s_entries_Freg_Tcmp[8][4] , \s_entries_Freg_Tcmp[8][3] , 
        \s_entries_Freg_Tcmp[8][2] , \s_entries_Freg_Tcmp[8][1] , 
        \s_entries_Freg_Tcmp[8][0] }) );
  NRegister_N32_98 EntrReg_i_9 ( .clk(BTB_clk), .reset(n332), .data_in({n219, 
        n216, n213, n210, n207, n204, n201, n198, n195, n192, n189, n186, n183, 
        n180, n177, n174, n171, n168, n165, n162, n159, n156, n153, n150, n147, 
        n144, n141, n138, n135, n132, n129, n126}), .enable(n17), .load(
        s_regenabl_entry[22]), .data_out({\s_entries_Freg_Tcmp[9][31] , 
        \s_entries_Freg_Tcmp[9][30] , \s_entries_Freg_Tcmp[9][29] , 
        \s_entries_Freg_Tcmp[9][28] , \s_entries_Freg_Tcmp[9][27] , 
        \s_entries_Freg_Tcmp[9][26] , \s_entries_Freg_Tcmp[9][25] , 
        \s_entries_Freg_Tcmp[9][24] , \s_entries_Freg_Tcmp[9][23] , 
        \s_entries_Freg_Tcmp[9][22] , \s_entries_Freg_Tcmp[9][21] , 
        \s_entries_Freg_Tcmp[9][20] , \s_entries_Freg_Tcmp[9][19] , 
        \s_entries_Freg_Tcmp[9][18] , \s_entries_Freg_Tcmp[9][17] , 
        \s_entries_Freg_Tcmp[9][16] , \s_entries_Freg_Tcmp[9][15] , 
        \s_entries_Freg_Tcmp[9][14] , \s_entries_Freg_Tcmp[9][13] , 
        \s_entries_Freg_Tcmp[9][12] , \s_entries_Freg_Tcmp[9][11] , 
        \s_entries_Freg_Tcmp[9][10] , \s_entries_Freg_Tcmp[9][9] , 
        \s_entries_Freg_Tcmp[9][8] , \s_entries_Freg_Tcmp[9][7] , 
        \s_entries_Freg_Tcmp[9][6] , \s_entries_Freg_Tcmp[9][5] , 
        \s_entries_Freg_Tcmp[9][4] , \s_entries_Freg_Tcmp[9][3] , 
        \s_entries_Freg_Tcmp[9][2] , \s_entries_Freg_Tcmp[9][1] , 
        \s_entries_Freg_Tcmp[9][0] }) );
  NRegister_N32_97 EntrReg_i_10 ( .clk(BTB_clk), .reset(n332), .data_in({n219, 
        n216, n213, n210, n207, n204, n201, n198, n195, n192, n189, n186, n183, 
        n180, n177, n174, n171, n168, n165, n162, n159, n156, n153, n150, n147, 
        n144, n141, n138, n135, n132, n129, n126}), .enable(n17), .load(
        s_regenabl_entry[21]), .data_out({\s_entries_Freg_Tcmp[10][31] , 
        \s_entries_Freg_Tcmp[10][30] , \s_entries_Freg_Tcmp[10][29] , 
        \s_entries_Freg_Tcmp[10][28] , \s_entries_Freg_Tcmp[10][27] , 
        \s_entries_Freg_Tcmp[10][26] , \s_entries_Freg_Tcmp[10][25] , 
        \s_entries_Freg_Tcmp[10][24] , \s_entries_Freg_Tcmp[10][23] , 
        \s_entries_Freg_Tcmp[10][22] , \s_entries_Freg_Tcmp[10][21] , 
        \s_entries_Freg_Tcmp[10][20] , \s_entries_Freg_Tcmp[10][19] , 
        \s_entries_Freg_Tcmp[10][18] , \s_entries_Freg_Tcmp[10][17] , 
        \s_entries_Freg_Tcmp[10][16] , \s_entries_Freg_Tcmp[10][15] , 
        \s_entries_Freg_Tcmp[10][14] , \s_entries_Freg_Tcmp[10][13] , 
        \s_entries_Freg_Tcmp[10][12] , \s_entries_Freg_Tcmp[10][11] , 
        \s_entries_Freg_Tcmp[10][10] , \s_entries_Freg_Tcmp[10][9] , 
        \s_entries_Freg_Tcmp[10][8] , \s_entries_Freg_Tcmp[10][7] , 
        \s_entries_Freg_Tcmp[10][6] , \s_entries_Freg_Tcmp[10][5] , 
        \s_entries_Freg_Tcmp[10][4] , \s_entries_Freg_Tcmp[10][3] , 
        \s_entries_Freg_Tcmp[10][2] , \s_entries_Freg_Tcmp[10][1] , 
        \s_entries_Freg_Tcmp[10][0] }) );
  NRegister_N32_96 EntrReg_i_11 ( .clk(BTB_clk), .reset(n332), .data_in({n219, 
        n216, n213, n210, n207, n204, n201, n198, n195, n192, n189, n186, n183, 
        n180, n177, n174, n171, n168, n165, n162, n159, n156, n153, n150, n147, 
        n144, n141, n138, n135, n132, n129, n126}), .enable(n17), .load(
        s_regenabl_entry[20]), .data_out({\s_entries_Freg_Tcmp[11][31] , 
        \s_entries_Freg_Tcmp[11][30] , \s_entries_Freg_Tcmp[11][29] , 
        \s_entries_Freg_Tcmp[11][28] , \s_entries_Freg_Tcmp[11][27] , 
        \s_entries_Freg_Tcmp[11][26] , \s_entries_Freg_Tcmp[11][25] , 
        \s_entries_Freg_Tcmp[11][24] , \s_entries_Freg_Tcmp[11][23] , 
        \s_entries_Freg_Tcmp[11][22] , \s_entries_Freg_Tcmp[11][21] , 
        \s_entries_Freg_Tcmp[11][20] , \s_entries_Freg_Tcmp[11][19] , 
        \s_entries_Freg_Tcmp[11][18] , \s_entries_Freg_Tcmp[11][17] , 
        \s_entries_Freg_Tcmp[11][16] , \s_entries_Freg_Tcmp[11][15] , 
        \s_entries_Freg_Tcmp[11][14] , \s_entries_Freg_Tcmp[11][13] , 
        \s_entries_Freg_Tcmp[11][12] , \s_entries_Freg_Tcmp[11][11] , 
        \s_entries_Freg_Tcmp[11][10] , \s_entries_Freg_Tcmp[11][9] , 
        \s_entries_Freg_Tcmp[11][8] , \s_entries_Freg_Tcmp[11][7] , 
        \s_entries_Freg_Tcmp[11][6] , \s_entries_Freg_Tcmp[11][5] , 
        \s_entries_Freg_Tcmp[11][4] , \s_entries_Freg_Tcmp[11][3] , 
        \s_entries_Freg_Tcmp[11][2] , \s_entries_Freg_Tcmp[11][1] , 
        \s_entries_Freg_Tcmp[11][0] }) );
  NRegister_N32_95 EntrReg_i_12 ( .clk(BTB_clk), .reset(n332), .data_in({n220, 
        n217, n214, n211, n208, n205, n202, n199, n196, n193, n190, n187, n184, 
        n181, n178, n175, n172, n169, n166, n163, n160, n157, n154, n151, n148, 
        n145, n142, n139, n136, n133, n130, n127}), .enable(n18), .load(
        s_regenabl_entry[19]), .data_out({\s_entries_Freg_Tcmp[12][31] , 
        \s_entries_Freg_Tcmp[12][30] , \s_entries_Freg_Tcmp[12][29] , 
        \s_entries_Freg_Tcmp[12][28] , \s_entries_Freg_Tcmp[12][27] , 
        \s_entries_Freg_Tcmp[12][26] , \s_entries_Freg_Tcmp[12][25] , 
        \s_entries_Freg_Tcmp[12][24] , \s_entries_Freg_Tcmp[12][23] , 
        \s_entries_Freg_Tcmp[12][22] , \s_entries_Freg_Tcmp[12][21] , 
        \s_entries_Freg_Tcmp[12][20] , \s_entries_Freg_Tcmp[12][19] , 
        \s_entries_Freg_Tcmp[12][18] , \s_entries_Freg_Tcmp[12][17] , 
        \s_entries_Freg_Tcmp[12][16] , \s_entries_Freg_Tcmp[12][15] , 
        \s_entries_Freg_Tcmp[12][14] , \s_entries_Freg_Tcmp[12][13] , 
        \s_entries_Freg_Tcmp[12][12] , \s_entries_Freg_Tcmp[12][11] , 
        \s_entries_Freg_Tcmp[12][10] , \s_entries_Freg_Tcmp[12][9] , 
        \s_entries_Freg_Tcmp[12][8] , \s_entries_Freg_Tcmp[12][7] , 
        \s_entries_Freg_Tcmp[12][6] , \s_entries_Freg_Tcmp[12][5] , 
        \s_entries_Freg_Tcmp[12][4] , \s_entries_Freg_Tcmp[12][3] , 
        \s_entries_Freg_Tcmp[12][2] , \s_entries_Freg_Tcmp[12][1] , 
        \s_entries_Freg_Tcmp[12][0] }) );
  NRegister_N32_94 EntrReg_i_13 ( .clk(BTB_clk), .reset(n332), .data_in({n220, 
        n217, n214, n211, n208, n205, n202, n199, n196, n193, n190, n187, n184, 
        n181, n178, n175, n172, n169, n166, n163, n160, n157, n154, n151, n148, 
        n145, n142, n139, n136, n133, n130, n127}), .enable(n18), .load(
        s_regenabl_entry[18]), .data_out({\s_entries_Freg_Tcmp[13][31] , 
        \s_entries_Freg_Tcmp[13][30] , \s_entries_Freg_Tcmp[13][29] , 
        \s_entries_Freg_Tcmp[13][28] , \s_entries_Freg_Tcmp[13][27] , 
        \s_entries_Freg_Tcmp[13][26] , \s_entries_Freg_Tcmp[13][25] , 
        \s_entries_Freg_Tcmp[13][24] , \s_entries_Freg_Tcmp[13][23] , 
        \s_entries_Freg_Tcmp[13][22] , \s_entries_Freg_Tcmp[13][21] , 
        \s_entries_Freg_Tcmp[13][20] , \s_entries_Freg_Tcmp[13][19] , 
        \s_entries_Freg_Tcmp[13][18] , \s_entries_Freg_Tcmp[13][17] , 
        \s_entries_Freg_Tcmp[13][16] , \s_entries_Freg_Tcmp[13][15] , 
        \s_entries_Freg_Tcmp[13][14] , \s_entries_Freg_Tcmp[13][13] , 
        \s_entries_Freg_Tcmp[13][12] , \s_entries_Freg_Tcmp[13][11] , 
        \s_entries_Freg_Tcmp[13][10] , \s_entries_Freg_Tcmp[13][9] , 
        \s_entries_Freg_Tcmp[13][8] , \s_entries_Freg_Tcmp[13][7] , 
        \s_entries_Freg_Tcmp[13][6] , \s_entries_Freg_Tcmp[13][5] , 
        \s_entries_Freg_Tcmp[13][4] , \s_entries_Freg_Tcmp[13][3] , 
        \s_entries_Freg_Tcmp[13][2] , \s_entries_Freg_Tcmp[13][1] , 
        \s_entries_Freg_Tcmp[13][0] }) );
  NRegister_N32_93 EntrReg_i_14 ( .clk(BTB_clk), .reset(n332), .data_in({n220, 
        n217, n214, n211, n208, n205, n202, n199, n196, n193, n190, n187, n184, 
        n181, n178, n175, n172, n169, n166, n163, n160, n157, n154, n151, n148, 
        n145, n142, n139, n136, n133, n130, n127}), .enable(n18), .load(
        s_regenabl_entry[17]), .data_out({\s_entries_Freg_Tcmp[14][31] , 
        \s_entries_Freg_Tcmp[14][30] , \s_entries_Freg_Tcmp[14][29] , 
        \s_entries_Freg_Tcmp[14][28] , \s_entries_Freg_Tcmp[14][27] , 
        \s_entries_Freg_Tcmp[14][26] , \s_entries_Freg_Tcmp[14][25] , 
        \s_entries_Freg_Tcmp[14][24] , \s_entries_Freg_Tcmp[14][23] , 
        \s_entries_Freg_Tcmp[14][22] , \s_entries_Freg_Tcmp[14][21] , 
        \s_entries_Freg_Tcmp[14][20] , \s_entries_Freg_Tcmp[14][19] , 
        \s_entries_Freg_Tcmp[14][18] , \s_entries_Freg_Tcmp[14][17] , 
        \s_entries_Freg_Tcmp[14][16] , \s_entries_Freg_Tcmp[14][15] , 
        \s_entries_Freg_Tcmp[14][14] , \s_entries_Freg_Tcmp[14][13] , 
        \s_entries_Freg_Tcmp[14][12] , \s_entries_Freg_Tcmp[14][11] , 
        \s_entries_Freg_Tcmp[14][10] , \s_entries_Freg_Tcmp[14][9] , 
        \s_entries_Freg_Tcmp[14][8] , \s_entries_Freg_Tcmp[14][7] , 
        \s_entries_Freg_Tcmp[14][6] , \s_entries_Freg_Tcmp[14][5] , 
        \s_entries_Freg_Tcmp[14][4] , \s_entries_Freg_Tcmp[14][3] , 
        \s_entries_Freg_Tcmp[14][2] , \s_entries_Freg_Tcmp[14][1] , 
        \s_entries_Freg_Tcmp[14][0] }) );
  NRegister_N32_92 EntrReg_i_15 ( .clk(BTB_clk), .reset(n332), .data_in({n220, 
        n217, n214, n211, n208, n205, n202, n199, n196, n193, n190, n187, n184, 
        n181, n178, n175, n172, n169, n166, n163, n160, n157, n154, n151, n148, 
        n145, n142, n139, n136, n133, n130, n127}), .enable(n18), .load(
        s_regenabl_entry[16]), .data_out({\s_entries_Freg_Tcmp[15][31] , 
        \s_entries_Freg_Tcmp[15][30] , \s_entries_Freg_Tcmp[15][29] , 
        \s_entries_Freg_Tcmp[15][28] , \s_entries_Freg_Tcmp[15][27] , 
        \s_entries_Freg_Tcmp[15][26] , \s_entries_Freg_Tcmp[15][25] , 
        \s_entries_Freg_Tcmp[15][24] , \s_entries_Freg_Tcmp[15][23] , 
        \s_entries_Freg_Tcmp[15][22] , \s_entries_Freg_Tcmp[15][21] , 
        \s_entries_Freg_Tcmp[15][20] , \s_entries_Freg_Tcmp[15][19] , 
        \s_entries_Freg_Tcmp[15][18] , \s_entries_Freg_Tcmp[15][17] , 
        \s_entries_Freg_Tcmp[15][16] , \s_entries_Freg_Tcmp[15][15] , 
        \s_entries_Freg_Tcmp[15][14] , \s_entries_Freg_Tcmp[15][13] , 
        \s_entries_Freg_Tcmp[15][12] , \s_entries_Freg_Tcmp[15][11] , 
        \s_entries_Freg_Tcmp[15][10] , \s_entries_Freg_Tcmp[15][9] , 
        \s_entries_Freg_Tcmp[15][8] , \s_entries_Freg_Tcmp[15][7] , 
        \s_entries_Freg_Tcmp[15][6] , \s_entries_Freg_Tcmp[15][5] , 
        \s_entries_Freg_Tcmp[15][4] , \s_entries_Freg_Tcmp[15][3] , 
        \s_entries_Freg_Tcmp[15][2] , \s_entries_Freg_Tcmp[15][1] , 
        \s_entries_Freg_Tcmp[15][0] }) );
  NRegister_N32_91 EntrReg_i_16 ( .clk(BTB_clk), .reset(n332), .data_in({n220, 
        n217, n214, n211, n208, n205, n202, n199, n196, n193, n190, n187, n184, 
        n181, n178, n175, n172, n169, n166, n163, n160, n157, n154, n151, n148, 
        n145, n142, n139, n136, n133, n130, n127}), .enable(n18), .load(
        s_regenabl_entry[15]), .data_out({\s_entries_Freg_Tcmp[16][31] , 
        \s_entries_Freg_Tcmp[16][30] , \s_entries_Freg_Tcmp[16][29] , 
        \s_entries_Freg_Tcmp[16][28] , \s_entries_Freg_Tcmp[16][27] , 
        \s_entries_Freg_Tcmp[16][26] , \s_entries_Freg_Tcmp[16][25] , 
        \s_entries_Freg_Tcmp[16][24] , \s_entries_Freg_Tcmp[16][23] , 
        \s_entries_Freg_Tcmp[16][22] , \s_entries_Freg_Tcmp[16][21] , 
        \s_entries_Freg_Tcmp[16][20] , \s_entries_Freg_Tcmp[16][19] , 
        \s_entries_Freg_Tcmp[16][18] , \s_entries_Freg_Tcmp[16][17] , 
        \s_entries_Freg_Tcmp[16][16] , \s_entries_Freg_Tcmp[16][15] , 
        \s_entries_Freg_Tcmp[16][14] , \s_entries_Freg_Tcmp[16][13] , 
        \s_entries_Freg_Tcmp[16][12] , \s_entries_Freg_Tcmp[16][11] , 
        \s_entries_Freg_Tcmp[16][10] , \s_entries_Freg_Tcmp[16][9] , 
        \s_entries_Freg_Tcmp[16][8] , \s_entries_Freg_Tcmp[16][7] , 
        \s_entries_Freg_Tcmp[16][6] , \s_entries_Freg_Tcmp[16][5] , 
        \s_entries_Freg_Tcmp[16][4] , \s_entries_Freg_Tcmp[16][3] , 
        \s_entries_Freg_Tcmp[16][2] , \s_entries_Freg_Tcmp[16][1] , 
        \s_entries_Freg_Tcmp[16][0] }) );
  NRegister_N32_90 EntrReg_i_17 ( .clk(BTB_clk), .reset(n331), .data_in({n220, 
        n217, n214, n211, n208, n205, n202, n199, n196, n193, n190, n187, n184, 
        n181, n178, n175, n172, n169, n166, n163, n160, n157, n154, n151, n148, 
        n145, n142, n139, n136, n133, n130, n127}), .enable(n18), .load(
        s_regenabl_entry[14]), .data_out({\s_entries_Freg_Tcmp[17][31] , 
        \s_entries_Freg_Tcmp[17][30] , \s_entries_Freg_Tcmp[17][29] , 
        \s_entries_Freg_Tcmp[17][28] , \s_entries_Freg_Tcmp[17][27] , 
        \s_entries_Freg_Tcmp[17][26] , \s_entries_Freg_Tcmp[17][25] , 
        \s_entries_Freg_Tcmp[17][24] , \s_entries_Freg_Tcmp[17][23] , 
        \s_entries_Freg_Tcmp[17][22] , \s_entries_Freg_Tcmp[17][21] , 
        \s_entries_Freg_Tcmp[17][20] , \s_entries_Freg_Tcmp[17][19] , 
        \s_entries_Freg_Tcmp[17][18] , \s_entries_Freg_Tcmp[17][17] , 
        \s_entries_Freg_Tcmp[17][16] , \s_entries_Freg_Tcmp[17][15] , 
        \s_entries_Freg_Tcmp[17][14] , \s_entries_Freg_Tcmp[17][13] , 
        \s_entries_Freg_Tcmp[17][12] , \s_entries_Freg_Tcmp[17][11] , 
        \s_entries_Freg_Tcmp[17][10] , \s_entries_Freg_Tcmp[17][9] , 
        \s_entries_Freg_Tcmp[17][8] , \s_entries_Freg_Tcmp[17][7] , 
        \s_entries_Freg_Tcmp[17][6] , \s_entries_Freg_Tcmp[17][5] , 
        \s_entries_Freg_Tcmp[17][4] , \s_entries_Freg_Tcmp[17][3] , 
        \s_entries_Freg_Tcmp[17][2] , \s_entries_Freg_Tcmp[17][1] , 
        \s_entries_Freg_Tcmp[17][0] }) );
  NRegister_N32_89 EntrReg_i_18 ( .clk(BTB_clk), .reset(n331), .data_in({n220, 
        n217, n214, n211, n208, n205, n202, n199, n196, n193, n190, n187, n184, 
        n181, n178, n175, n172, n169, n166, n163, n160, n157, n154, n151, n148, 
        n145, n142, n139, n136, n133, n130, n127}), .enable(n18), .load(
        s_regenabl_entry[13]), .data_out({\s_entries_Freg_Tcmp[18][31] , 
        \s_entries_Freg_Tcmp[18][30] , \s_entries_Freg_Tcmp[18][29] , 
        \s_entries_Freg_Tcmp[18][28] , \s_entries_Freg_Tcmp[18][27] , 
        \s_entries_Freg_Tcmp[18][26] , \s_entries_Freg_Tcmp[18][25] , 
        \s_entries_Freg_Tcmp[18][24] , \s_entries_Freg_Tcmp[18][23] , 
        \s_entries_Freg_Tcmp[18][22] , \s_entries_Freg_Tcmp[18][21] , 
        \s_entries_Freg_Tcmp[18][20] , \s_entries_Freg_Tcmp[18][19] , 
        \s_entries_Freg_Tcmp[18][18] , \s_entries_Freg_Tcmp[18][17] , 
        \s_entries_Freg_Tcmp[18][16] , \s_entries_Freg_Tcmp[18][15] , 
        \s_entries_Freg_Tcmp[18][14] , \s_entries_Freg_Tcmp[18][13] , 
        \s_entries_Freg_Tcmp[18][12] , \s_entries_Freg_Tcmp[18][11] , 
        \s_entries_Freg_Tcmp[18][10] , \s_entries_Freg_Tcmp[18][9] , 
        \s_entries_Freg_Tcmp[18][8] , \s_entries_Freg_Tcmp[18][7] , 
        \s_entries_Freg_Tcmp[18][6] , \s_entries_Freg_Tcmp[18][5] , 
        \s_entries_Freg_Tcmp[18][4] , \s_entries_Freg_Tcmp[18][3] , 
        \s_entries_Freg_Tcmp[18][2] , \s_entries_Freg_Tcmp[18][1] , 
        \s_entries_Freg_Tcmp[18][0] }) );
  NRegister_N32_88 EntrReg_i_19 ( .clk(BTB_clk), .reset(n331), .data_in({n220, 
        n217, n214, n211, n208, n205, n202, n199, n196, n193, n190, n187, n184, 
        n181, n178, n175, n172, n169, n166, n163, n160, n157, n154, n151, n148, 
        n145, n142, n139, n136, n133, n130, n127}), .enable(n18), .load(
        s_regenabl_entry[12]), .data_out({\s_entries_Freg_Tcmp[19][31] , 
        \s_entries_Freg_Tcmp[19][30] , \s_entries_Freg_Tcmp[19][29] , 
        \s_entries_Freg_Tcmp[19][28] , \s_entries_Freg_Tcmp[19][27] , 
        \s_entries_Freg_Tcmp[19][26] , \s_entries_Freg_Tcmp[19][25] , 
        \s_entries_Freg_Tcmp[19][24] , \s_entries_Freg_Tcmp[19][23] , 
        \s_entries_Freg_Tcmp[19][22] , \s_entries_Freg_Tcmp[19][21] , 
        \s_entries_Freg_Tcmp[19][20] , \s_entries_Freg_Tcmp[19][19] , 
        \s_entries_Freg_Tcmp[19][18] , \s_entries_Freg_Tcmp[19][17] , 
        \s_entries_Freg_Tcmp[19][16] , \s_entries_Freg_Tcmp[19][15] , 
        \s_entries_Freg_Tcmp[19][14] , \s_entries_Freg_Tcmp[19][13] , 
        \s_entries_Freg_Tcmp[19][12] , \s_entries_Freg_Tcmp[19][11] , 
        \s_entries_Freg_Tcmp[19][10] , \s_entries_Freg_Tcmp[19][9] , 
        \s_entries_Freg_Tcmp[19][8] , \s_entries_Freg_Tcmp[19][7] , 
        \s_entries_Freg_Tcmp[19][6] , \s_entries_Freg_Tcmp[19][5] , 
        \s_entries_Freg_Tcmp[19][4] , \s_entries_Freg_Tcmp[19][3] , 
        \s_entries_Freg_Tcmp[19][2] , \s_entries_Freg_Tcmp[19][1] , 
        \s_entries_Freg_Tcmp[19][0] }) );
  NRegister_N32_87 EntrReg_i_20 ( .clk(BTB_clk), .reset(n331), .data_in({n220, 
        n217, n214, n211, n208, n205, n202, n199, n196, n193, n190, n187, n184, 
        n181, n178, n175, n172, n169, n166, n163, n160, n157, n154, n151, n148, 
        n145, n142, n139, n136, n133, n130, n127}), .enable(n18), .load(
        s_regenabl_entry[11]), .data_out({\s_entries_Freg_Tcmp[20][31] , 
        \s_entries_Freg_Tcmp[20][30] , \s_entries_Freg_Tcmp[20][29] , 
        \s_entries_Freg_Tcmp[20][28] , \s_entries_Freg_Tcmp[20][27] , 
        \s_entries_Freg_Tcmp[20][26] , \s_entries_Freg_Tcmp[20][25] , 
        \s_entries_Freg_Tcmp[20][24] , \s_entries_Freg_Tcmp[20][23] , 
        \s_entries_Freg_Tcmp[20][22] , \s_entries_Freg_Tcmp[20][21] , 
        \s_entries_Freg_Tcmp[20][20] , \s_entries_Freg_Tcmp[20][19] , 
        \s_entries_Freg_Tcmp[20][18] , \s_entries_Freg_Tcmp[20][17] , 
        \s_entries_Freg_Tcmp[20][16] , \s_entries_Freg_Tcmp[20][15] , 
        \s_entries_Freg_Tcmp[20][14] , \s_entries_Freg_Tcmp[20][13] , 
        \s_entries_Freg_Tcmp[20][12] , \s_entries_Freg_Tcmp[20][11] , 
        \s_entries_Freg_Tcmp[20][10] , \s_entries_Freg_Tcmp[20][9] , 
        \s_entries_Freg_Tcmp[20][8] , \s_entries_Freg_Tcmp[20][7] , 
        \s_entries_Freg_Tcmp[20][6] , \s_entries_Freg_Tcmp[20][5] , 
        \s_entries_Freg_Tcmp[20][4] , \s_entries_Freg_Tcmp[20][3] , 
        \s_entries_Freg_Tcmp[20][2] , \s_entries_Freg_Tcmp[20][1] , 
        \s_entries_Freg_Tcmp[20][0] }) );
  NRegister_N32_86 EntrReg_i_21 ( .clk(BTB_clk), .reset(n331), .data_in({n220, 
        n217, n214, n211, n208, n205, n202, n199, n196, n193, n190, n187, n184, 
        n181, n178, n175, n172, n169, n166, n163, n160, n157, n154, n151, n148, 
        n145, n142, n139, n136, n133, n130, n127}), .enable(n18), .load(
        s_regenabl_entry[10]), .data_out({\s_entries_Freg_Tcmp[21][31] , 
        \s_entries_Freg_Tcmp[21][30] , \s_entries_Freg_Tcmp[21][29] , 
        \s_entries_Freg_Tcmp[21][28] , \s_entries_Freg_Tcmp[21][27] , 
        \s_entries_Freg_Tcmp[21][26] , \s_entries_Freg_Tcmp[21][25] , 
        \s_entries_Freg_Tcmp[21][24] , \s_entries_Freg_Tcmp[21][23] , 
        \s_entries_Freg_Tcmp[21][22] , \s_entries_Freg_Tcmp[21][21] , 
        \s_entries_Freg_Tcmp[21][20] , \s_entries_Freg_Tcmp[21][19] , 
        \s_entries_Freg_Tcmp[21][18] , \s_entries_Freg_Tcmp[21][17] , 
        \s_entries_Freg_Tcmp[21][16] , \s_entries_Freg_Tcmp[21][15] , 
        \s_entries_Freg_Tcmp[21][14] , \s_entries_Freg_Tcmp[21][13] , 
        \s_entries_Freg_Tcmp[21][12] , \s_entries_Freg_Tcmp[21][11] , 
        \s_entries_Freg_Tcmp[21][10] , \s_entries_Freg_Tcmp[21][9] , 
        \s_entries_Freg_Tcmp[21][8] , \s_entries_Freg_Tcmp[21][7] , 
        \s_entries_Freg_Tcmp[21][6] , \s_entries_Freg_Tcmp[21][5] , 
        \s_entries_Freg_Tcmp[21][4] , \s_entries_Freg_Tcmp[21][3] , 
        \s_entries_Freg_Tcmp[21][2] , \s_entries_Freg_Tcmp[21][1] , 
        \s_entries_Freg_Tcmp[21][0] }) );
  NRegister_N32_85 EntrReg_i_22 ( .clk(BTB_clk), .reset(n331), .data_in({n220, 
        n217, n214, n211, n208, n205, n202, n199, n196, n193, n190, n187, n184, 
        n181, n178, n175, n172, n169, n166, n163, n160, n157, n154, n151, n148, 
        n145, n142, n139, n136, n133, n130, n127}), .enable(n18), .load(
        s_regenabl_entry[9]), .data_out({\s_entries_Freg_Tcmp[22][31] , 
        \s_entries_Freg_Tcmp[22][30] , \s_entries_Freg_Tcmp[22][29] , 
        \s_entries_Freg_Tcmp[22][28] , \s_entries_Freg_Tcmp[22][27] , 
        \s_entries_Freg_Tcmp[22][26] , \s_entries_Freg_Tcmp[22][25] , 
        \s_entries_Freg_Tcmp[22][24] , \s_entries_Freg_Tcmp[22][23] , 
        \s_entries_Freg_Tcmp[22][22] , \s_entries_Freg_Tcmp[22][21] , 
        \s_entries_Freg_Tcmp[22][20] , \s_entries_Freg_Tcmp[22][19] , 
        \s_entries_Freg_Tcmp[22][18] , \s_entries_Freg_Tcmp[22][17] , 
        \s_entries_Freg_Tcmp[22][16] , \s_entries_Freg_Tcmp[22][15] , 
        \s_entries_Freg_Tcmp[22][14] , \s_entries_Freg_Tcmp[22][13] , 
        \s_entries_Freg_Tcmp[22][12] , \s_entries_Freg_Tcmp[22][11] , 
        \s_entries_Freg_Tcmp[22][10] , \s_entries_Freg_Tcmp[22][9] , 
        \s_entries_Freg_Tcmp[22][8] , \s_entries_Freg_Tcmp[22][7] , 
        \s_entries_Freg_Tcmp[22][6] , \s_entries_Freg_Tcmp[22][5] , 
        \s_entries_Freg_Tcmp[22][4] , \s_entries_Freg_Tcmp[22][3] , 
        \s_entries_Freg_Tcmp[22][2] , \s_entries_Freg_Tcmp[22][1] , 
        \s_entries_Freg_Tcmp[22][0] }) );
  NRegister_N32_84 EntrReg_i_23 ( .clk(BTB_clk), .reset(n331), .data_in({n220, 
        n217, n214, n211, n208, n205, n202, n199, n196, n193, n190, n187, n184, 
        n181, n178, n175, n172, n169, n166, n163, n160, n157, n154, n151, n148, 
        n145, n142, n139, n136, n133, n130, n127}), .enable(n18), .load(
        s_regenabl_entry[8]), .data_out({\s_entries_Freg_Tcmp[23][31] , 
        \s_entries_Freg_Tcmp[23][30] , \s_entries_Freg_Tcmp[23][29] , 
        \s_entries_Freg_Tcmp[23][28] , \s_entries_Freg_Tcmp[23][27] , 
        \s_entries_Freg_Tcmp[23][26] , \s_entries_Freg_Tcmp[23][25] , 
        \s_entries_Freg_Tcmp[23][24] , \s_entries_Freg_Tcmp[23][23] , 
        \s_entries_Freg_Tcmp[23][22] , \s_entries_Freg_Tcmp[23][21] , 
        \s_entries_Freg_Tcmp[23][20] , \s_entries_Freg_Tcmp[23][19] , 
        \s_entries_Freg_Tcmp[23][18] , \s_entries_Freg_Tcmp[23][17] , 
        \s_entries_Freg_Tcmp[23][16] , \s_entries_Freg_Tcmp[23][15] , 
        \s_entries_Freg_Tcmp[23][14] , \s_entries_Freg_Tcmp[23][13] , 
        \s_entries_Freg_Tcmp[23][12] , \s_entries_Freg_Tcmp[23][11] , 
        \s_entries_Freg_Tcmp[23][10] , \s_entries_Freg_Tcmp[23][9] , 
        \s_entries_Freg_Tcmp[23][8] , \s_entries_Freg_Tcmp[23][7] , 
        \s_entries_Freg_Tcmp[23][6] , \s_entries_Freg_Tcmp[23][5] , 
        \s_entries_Freg_Tcmp[23][4] , \s_entries_Freg_Tcmp[23][3] , 
        \s_entries_Freg_Tcmp[23][2] , \s_entries_Freg_Tcmp[23][1] , 
        \s_entries_Freg_Tcmp[23][0] }) );
  NRegister_N32_83 EntrReg_i_24 ( .clk(BTB_clk), .reset(n331), .data_in({n221, 
        n218, n215, n212, n209, n206, n203, n200, n197, n194, n191, n188, n185, 
        n182, n179, n176, n173, n170, n167, n164, n161, n158, n155, n152, n149, 
        n146, n143, n140, n137, n134, n131, n128}), .enable(n19), .load(
        s_regenabl_entry[7]), .data_out({\s_entries_Freg_Tcmp[24][31] , 
        \s_entries_Freg_Tcmp[24][30] , \s_entries_Freg_Tcmp[24][29] , 
        \s_entries_Freg_Tcmp[24][28] , \s_entries_Freg_Tcmp[24][27] , 
        \s_entries_Freg_Tcmp[24][26] , \s_entries_Freg_Tcmp[24][25] , 
        \s_entries_Freg_Tcmp[24][24] , \s_entries_Freg_Tcmp[24][23] , 
        \s_entries_Freg_Tcmp[24][22] , \s_entries_Freg_Tcmp[24][21] , 
        \s_entries_Freg_Tcmp[24][20] , \s_entries_Freg_Tcmp[24][19] , 
        \s_entries_Freg_Tcmp[24][18] , \s_entries_Freg_Tcmp[24][17] , 
        \s_entries_Freg_Tcmp[24][16] , \s_entries_Freg_Tcmp[24][15] , 
        \s_entries_Freg_Tcmp[24][14] , \s_entries_Freg_Tcmp[24][13] , 
        \s_entries_Freg_Tcmp[24][12] , \s_entries_Freg_Tcmp[24][11] , 
        \s_entries_Freg_Tcmp[24][10] , \s_entries_Freg_Tcmp[24][9] , 
        \s_entries_Freg_Tcmp[24][8] , \s_entries_Freg_Tcmp[24][7] , 
        \s_entries_Freg_Tcmp[24][6] , \s_entries_Freg_Tcmp[24][5] , 
        \s_entries_Freg_Tcmp[24][4] , \s_entries_Freg_Tcmp[24][3] , 
        \s_entries_Freg_Tcmp[24][2] , \s_entries_Freg_Tcmp[24][1] , 
        \s_entries_Freg_Tcmp[24][0] }) );
  NRegister_N32_82 EntrReg_i_25 ( .clk(BTB_clk), .reset(n331), .data_in({n221, 
        n218, n215, n212, n209, n206, n203, n200, n197, n194, n191, n188, n185, 
        n182, n179, n176, n173, n170, n167, n164, n161, n158, n155, n152, n149, 
        n146, n143, n140, n137, n134, n131, n128}), .enable(n19), .load(
        s_regenabl_entry[6]), .data_out({\s_entries_Freg_Tcmp[25][31] , 
        \s_entries_Freg_Tcmp[25][30] , \s_entries_Freg_Tcmp[25][29] , 
        \s_entries_Freg_Tcmp[25][28] , \s_entries_Freg_Tcmp[25][27] , 
        \s_entries_Freg_Tcmp[25][26] , \s_entries_Freg_Tcmp[25][25] , 
        \s_entries_Freg_Tcmp[25][24] , \s_entries_Freg_Tcmp[25][23] , 
        \s_entries_Freg_Tcmp[25][22] , \s_entries_Freg_Tcmp[25][21] , 
        \s_entries_Freg_Tcmp[25][20] , \s_entries_Freg_Tcmp[25][19] , 
        \s_entries_Freg_Tcmp[25][18] , \s_entries_Freg_Tcmp[25][17] , 
        \s_entries_Freg_Tcmp[25][16] , \s_entries_Freg_Tcmp[25][15] , 
        \s_entries_Freg_Tcmp[25][14] , \s_entries_Freg_Tcmp[25][13] , 
        \s_entries_Freg_Tcmp[25][12] , \s_entries_Freg_Tcmp[25][11] , 
        \s_entries_Freg_Tcmp[25][10] , \s_entries_Freg_Tcmp[25][9] , 
        \s_entries_Freg_Tcmp[25][8] , \s_entries_Freg_Tcmp[25][7] , 
        \s_entries_Freg_Tcmp[25][6] , \s_entries_Freg_Tcmp[25][5] , 
        \s_entries_Freg_Tcmp[25][4] , \s_entries_Freg_Tcmp[25][3] , 
        \s_entries_Freg_Tcmp[25][2] , \s_entries_Freg_Tcmp[25][1] , 
        \s_entries_Freg_Tcmp[25][0] }) );
  NRegister_N32_81 EntrReg_i_26 ( .clk(BTB_clk), .reset(n331), .data_in({n221, 
        n218, n215, n212, n209, n206, n203, n200, n197, n194, n191, n188, n185, 
        n182, n179, n176, n173, n170, n167, n164, n161, n158, n155, n152, n149, 
        n146, n143, n140, n137, n134, n131, n128}), .enable(n19), .load(
        s_regenabl_entry[5]), .data_out({\s_entries_Freg_Tcmp[26][31] , 
        \s_entries_Freg_Tcmp[26][30] , \s_entries_Freg_Tcmp[26][29] , 
        \s_entries_Freg_Tcmp[26][28] , \s_entries_Freg_Tcmp[26][27] , 
        \s_entries_Freg_Tcmp[26][26] , \s_entries_Freg_Tcmp[26][25] , 
        \s_entries_Freg_Tcmp[26][24] , \s_entries_Freg_Tcmp[26][23] , 
        \s_entries_Freg_Tcmp[26][22] , \s_entries_Freg_Tcmp[26][21] , 
        \s_entries_Freg_Tcmp[26][20] , \s_entries_Freg_Tcmp[26][19] , 
        \s_entries_Freg_Tcmp[26][18] , \s_entries_Freg_Tcmp[26][17] , 
        \s_entries_Freg_Tcmp[26][16] , \s_entries_Freg_Tcmp[26][15] , 
        \s_entries_Freg_Tcmp[26][14] , \s_entries_Freg_Tcmp[26][13] , 
        \s_entries_Freg_Tcmp[26][12] , \s_entries_Freg_Tcmp[26][11] , 
        \s_entries_Freg_Tcmp[26][10] , \s_entries_Freg_Tcmp[26][9] , 
        \s_entries_Freg_Tcmp[26][8] , \s_entries_Freg_Tcmp[26][7] , 
        \s_entries_Freg_Tcmp[26][6] , \s_entries_Freg_Tcmp[26][5] , 
        \s_entries_Freg_Tcmp[26][4] , \s_entries_Freg_Tcmp[26][3] , 
        \s_entries_Freg_Tcmp[26][2] , \s_entries_Freg_Tcmp[26][1] , 
        \s_entries_Freg_Tcmp[26][0] }) );
  NRegister_N32_80 EntrReg_i_27 ( .clk(BTB_clk), .reset(n331), .data_in({n221, 
        n218, n215, n212, n209, n206, n203, n200, n197, n194, n191, n188, n185, 
        n182, n179, n176, n173, n170, n167, n164, n161, n158, n155, n152, n149, 
        n146, n143, n140, n137, n134, n131, n128}), .enable(n19), .load(
        s_regenabl_entry[4]), .data_out({\s_entries_Freg_Tcmp[27][31] , 
        \s_entries_Freg_Tcmp[27][30] , \s_entries_Freg_Tcmp[27][29] , 
        \s_entries_Freg_Tcmp[27][28] , \s_entries_Freg_Tcmp[27][27] , 
        \s_entries_Freg_Tcmp[27][26] , \s_entries_Freg_Tcmp[27][25] , 
        \s_entries_Freg_Tcmp[27][24] , \s_entries_Freg_Tcmp[27][23] , 
        \s_entries_Freg_Tcmp[27][22] , \s_entries_Freg_Tcmp[27][21] , 
        \s_entries_Freg_Tcmp[27][20] , \s_entries_Freg_Tcmp[27][19] , 
        \s_entries_Freg_Tcmp[27][18] , \s_entries_Freg_Tcmp[27][17] , 
        \s_entries_Freg_Tcmp[27][16] , \s_entries_Freg_Tcmp[27][15] , 
        \s_entries_Freg_Tcmp[27][14] , \s_entries_Freg_Tcmp[27][13] , 
        \s_entries_Freg_Tcmp[27][12] , \s_entries_Freg_Tcmp[27][11] , 
        \s_entries_Freg_Tcmp[27][10] , \s_entries_Freg_Tcmp[27][9] , 
        \s_entries_Freg_Tcmp[27][8] , \s_entries_Freg_Tcmp[27][7] , 
        \s_entries_Freg_Tcmp[27][6] , \s_entries_Freg_Tcmp[27][5] , 
        \s_entries_Freg_Tcmp[27][4] , \s_entries_Freg_Tcmp[27][3] , 
        \s_entries_Freg_Tcmp[27][2] , \s_entries_Freg_Tcmp[27][1] , 
        \s_entries_Freg_Tcmp[27][0] }) );
  NRegister_N32_79 EntrReg_i_28 ( .clk(BTB_clk), .reset(n331), .data_in({n221, 
        n218, n215, n212, n209, n206, n203, n200, n197, n194, n191, n188, n185, 
        n182, n179, n176, n173, n170, n167, n164, n161, n158, n155, n152, n149, 
        n146, n143, n140, n137, n134, n131, n128}), .enable(n19), .load(
        s_regenabl_entry[3]), .data_out({\s_entries_Freg_Tcmp[28][31] , 
        \s_entries_Freg_Tcmp[28][30] , \s_entries_Freg_Tcmp[28][29] , 
        \s_entries_Freg_Tcmp[28][28] , \s_entries_Freg_Tcmp[28][27] , 
        \s_entries_Freg_Tcmp[28][26] , \s_entries_Freg_Tcmp[28][25] , 
        \s_entries_Freg_Tcmp[28][24] , \s_entries_Freg_Tcmp[28][23] , 
        \s_entries_Freg_Tcmp[28][22] , \s_entries_Freg_Tcmp[28][21] , 
        \s_entries_Freg_Tcmp[28][20] , \s_entries_Freg_Tcmp[28][19] , 
        \s_entries_Freg_Tcmp[28][18] , \s_entries_Freg_Tcmp[28][17] , 
        \s_entries_Freg_Tcmp[28][16] , \s_entries_Freg_Tcmp[28][15] , 
        \s_entries_Freg_Tcmp[28][14] , \s_entries_Freg_Tcmp[28][13] , 
        \s_entries_Freg_Tcmp[28][12] , \s_entries_Freg_Tcmp[28][11] , 
        \s_entries_Freg_Tcmp[28][10] , \s_entries_Freg_Tcmp[28][9] , 
        \s_entries_Freg_Tcmp[28][8] , \s_entries_Freg_Tcmp[28][7] , 
        \s_entries_Freg_Tcmp[28][6] , \s_entries_Freg_Tcmp[28][5] , 
        \s_entries_Freg_Tcmp[28][4] , \s_entries_Freg_Tcmp[28][3] , 
        \s_entries_Freg_Tcmp[28][2] , \s_entries_Freg_Tcmp[28][1] , 
        \s_entries_Freg_Tcmp[28][0] }) );
  NRegister_N32_78 EntrReg_i_29 ( .clk(BTB_clk), .reset(n330), .data_in({n221, 
        n218, n215, n212, n209, n206, n203, n200, n197, n194, n191, n188, n185, 
        n182, n179, n176, n173, n170, n167, n164, n161, n158, n155, n152, n149, 
        n146, n143, n140, n137, n134, n131, n128}), .enable(n19), .load(
        s_regenabl_entry[2]), .data_out({\s_entries_Freg_Tcmp[29][31] , 
        \s_entries_Freg_Tcmp[29][30] , \s_entries_Freg_Tcmp[29][29] , 
        \s_entries_Freg_Tcmp[29][28] , \s_entries_Freg_Tcmp[29][27] , 
        \s_entries_Freg_Tcmp[29][26] , \s_entries_Freg_Tcmp[29][25] , 
        \s_entries_Freg_Tcmp[29][24] , \s_entries_Freg_Tcmp[29][23] , 
        \s_entries_Freg_Tcmp[29][22] , \s_entries_Freg_Tcmp[29][21] , 
        \s_entries_Freg_Tcmp[29][20] , \s_entries_Freg_Tcmp[29][19] , 
        \s_entries_Freg_Tcmp[29][18] , \s_entries_Freg_Tcmp[29][17] , 
        \s_entries_Freg_Tcmp[29][16] , \s_entries_Freg_Tcmp[29][15] , 
        \s_entries_Freg_Tcmp[29][14] , \s_entries_Freg_Tcmp[29][13] , 
        \s_entries_Freg_Tcmp[29][12] , \s_entries_Freg_Tcmp[29][11] , 
        \s_entries_Freg_Tcmp[29][10] , \s_entries_Freg_Tcmp[29][9] , 
        \s_entries_Freg_Tcmp[29][8] , \s_entries_Freg_Tcmp[29][7] , 
        \s_entries_Freg_Tcmp[29][6] , \s_entries_Freg_Tcmp[29][5] , 
        \s_entries_Freg_Tcmp[29][4] , \s_entries_Freg_Tcmp[29][3] , 
        \s_entries_Freg_Tcmp[29][2] , \s_entries_Freg_Tcmp[29][1] , 
        \s_entries_Freg_Tcmp[29][0] }) );
  NRegister_N32_77 EntrReg_i_30 ( .clk(BTB_clk), .reset(n330), .data_in({n221, 
        n218, n215, n212, n209, n206, n203, n200, n197, n194, n191, n188, n185, 
        n182, n179, n176, n173, n170, n167, n164, n161, n158, n155, n152, n149, 
        n146, n143, n140, n137, n134, n131, n128}), .enable(n19), .load(
        s_regenabl_entry[1]), .data_out({\s_entries_Freg_Tcmp[30][31] , 
        \s_entries_Freg_Tcmp[30][30] , \s_entries_Freg_Tcmp[30][29] , 
        \s_entries_Freg_Tcmp[30][28] , \s_entries_Freg_Tcmp[30][27] , 
        \s_entries_Freg_Tcmp[30][26] , \s_entries_Freg_Tcmp[30][25] , 
        \s_entries_Freg_Tcmp[30][24] , \s_entries_Freg_Tcmp[30][23] , 
        \s_entries_Freg_Tcmp[30][22] , \s_entries_Freg_Tcmp[30][21] , 
        \s_entries_Freg_Tcmp[30][20] , \s_entries_Freg_Tcmp[30][19] , 
        \s_entries_Freg_Tcmp[30][18] , \s_entries_Freg_Tcmp[30][17] , 
        \s_entries_Freg_Tcmp[30][16] , \s_entries_Freg_Tcmp[30][15] , 
        \s_entries_Freg_Tcmp[30][14] , \s_entries_Freg_Tcmp[30][13] , 
        \s_entries_Freg_Tcmp[30][12] , \s_entries_Freg_Tcmp[30][11] , 
        \s_entries_Freg_Tcmp[30][10] , \s_entries_Freg_Tcmp[30][9] , 
        \s_entries_Freg_Tcmp[30][8] , \s_entries_Freg_Tcmp[30][7] , 
        \s_entries_Freg_Tcmp[30][6] , \s_entries_Freg_Tcmp[30][5] , 
        \s_entries_Freg_Tcmp[30][4] , \s_entries_Freg_Tcmp[30][3] , 
        \s_entries_Freg_Tcmp[30][2] , \s_entries_Freg_Tcmp[30][1] , 
        \s_entries_Freg_Tcmp[30][0] }) );
  NRegister_N32_76 EntrReg_i_31 ( .clk(BTB_clk), .reset(n330), .data_in({n221, 
        n218, n215, n212, n209, n206, n203, n200, n197, n194, n191, n188, n185, 
        n182, n179, n176, n173, n170, n167, n164, n161, n158, n155, n152, n149, 
        n146, n143, n140, n137, n134, n131, n128}), .enable(n19), .load(
        s_regenabl_entry[0]), .data_out({\s_entries_Freg_Tcmp[31][31] , 
        \s_entries_Freg_Tcmp[31][30] , \s_entries_Freg_Tcmp[31][29] , 
        \s_entries_Freg_Tcmp[31][28] , \s_entries_Freg_Tcmp[31][27] , 
        \s_entries_Freg_Tcmp[31][26] , \s_entries_Freg_Tcmp[31][25] , 
        \s_entries_Freg_Tcmp[31][24] , \s_entries_Freg_Tcmp[31][23] , 
        \s_entries_Freg_Tcmp[31][22] , \s_entries_Freg_Tcmp[31][21] , 
        \s_entries_Freg_Tcmp[31][20] , \s_entries_Freg_Tcmp[31][19] , 
        \s_entries_Freg_Tcmp[31][18] , \s_entries_Freg_Tcmp[31][17] , 
        \s_entries_Freg_Tcmp[31][16] , \s_entries_Freg_Tcmp[31][15] , 
        \s_entries_Freg_Tcmp[31][14] , \s_entries_Freg_Tcmp[31][13] , 
        \s_entries_Freg_Tcmp[31][12] , \s_entries_Freg_Tcmp[31][11] , 
        \s_entries_Freg_Tcmp[31][10] , \s_entries_Freg_Tcmp[31][9] , 
        \s_entries_Freg_Tcmp[31][8] , \s_entries_Freg_Tcmp[31][7] , 
        \s_entries_Freg_Tcmp[31][6] , \s_entries_Freg_Tcmp[31][5] , 
        \s_entries_Freg_Tcmp[31][4] , \s_entries_Freg_Tcmp[31][3] , 
        \s_entries_Freg_Tcmp[31][2] , \s_entries_Freg_Tcmp[31][1] , 
        \s_entries_Freg_Tcmp[31][0] }) );
  NRegister_N32_75 TargReg_i_0 ( .clk(BTB_clk), .reset(n330), .data_in({n125, 
        n120, n117, n114, n111, n108, n105, n102, n99, n96, n93, n90, n87, n84, 
        n81, n78, n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, 
        n39, n36, n33, n30}), .enable(n19), .load(s_regenabl_target[31]), 
        .data_out({\s_mux_signals[0][0][31] , \s_mux_signals[0][0][30] , 
        \s_mux_signals[0][0][29] , \s_mux_signals[0][0][28] , 
        \s_mux_signals[0][0][27] , \s_mux_signals[0][0][26] , 
        \s_mux_signals[0][0][25] , \s_mux_signals[0][0][24] , 
        \s_mux_signals[0][0][23] , \s_mux_signals[0][0][22] , 
        \s_mux_signals[0][0][21] , \s_mux_signals[0][0][20] , 
        \s_mux_signals[0][0][19] , \s_mux_signals[0][0][18] , 
        \s_mux_signals[0][0][17] , \s_mux_signals[0][0][16] , 
        \s_mux_signals[0][0][15] , \s_mux_signals[0][0][14] , 
        \s_mux_signals[0][0][13] , \s_mux_signals[0][0][12] , 
        \s_mux_signals[0][0][11] , \s_mux_signals[0][0][10] , 
        \s_mux_signals[0][0][9] , \s_mux_signals[0][0][8] , 
        \s_mux_signals[0][0][7] , \s_mux_signals[0][0][6] , 
        \s_mux_signals[0][0][5] , \s_mux_signals[0][0][4] , 
        \s_mux_signals[0][0][3] , \s_mux_signals[0][0][2] , 
        \s_mux_signals[0][0][1] , \s_mux_signals[0][0][0] }) );
  NRegister_N32_74 TargReg_i_1 ( .clk(BTB_clk), .reset(n330), .data_in({n125, 
        n120, n117, n114, n111, n108, n105, n102, n99, n96, n93, n90, n87, n84, 
        n81, n78, n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, 
        n39, n36, n33, n30}), .enable(n19), .load(s_regenabl_target[30]), 
        .data_out({\s_mux_signals[0][1][31] , \s_mux_signals[0][1][30] , 
        \s_mux_signals[0][1][29] , \s_mux_signals[0][1][28] , 
        \s_mux_signals[0][1][27] , \s_mux_signals[0][1][26] , 
        \s_mux_signals[0][1][25] , \s_mux_signals[0][1][24] , 
        \s_mux_signals[0][1][23] , \s_mux_signals[0][1][22] , 
        \s_mux_signals[0][1][21] , \s_mux_signals[0][1][20] , 
        \s_mux_signals[0][1][19] , \s_mux_signals[0][1][18] , 
        \s_mux_signals[0][1][17] , \s_mux_signals[0][1][16] , 
        \s_mux_signals[0][1][15] , \s_mux_signals[0][1][14] , 
        \s_mux_signals[0][1][13] , \s_mux_signals[0][1][12] , 
        \s_mux_signals[0][1][11] , \s_mux_signals[0][1][10] , 
        \s_mux_signals[0][1][9] , \s_mux_signals[0][1][8] , 
        \s_mux_signals[0][1][7] , \s_mux_signals[0][1][6] , 
        \s_mux_signals[0][1][5] , \s_mux_signals[0][1][4] , 
        \s_mux_signals[0][1][3] , \s_mux_signals[0][1][2] , 
        \s_mux_signals[0][1][1] , \s_mux_signals[0][1][0] }) );
  NRegister_N32_73 TargReg_i_2 ( .clk(BTB_clk), .reset(n330), .data_in({n124, 
        n120, n117, n114, n111, n108, n105, n102, n99, n96, n93, n90, n87, n84, 
        n81, n78, n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, 
        n39, n36, n33, n30}), .enable(n19), .load(s_regenabl_target[29]), 
        .data_out({\s_mux_signals[0][2][31] , \s_mux_signals[0][2][30] , 
        \s_mux_signals[0][2][29] , \s_mux_signals[0][2][28] , 
        \s_mux_signals[0][2][27] , \s_mux_signals[0][2][26] , 
        \s_mux_signals[0][2][25] , \s_mux_signals[0][2][24] , 
        \s_mux_signals[0][2][23] , \s_mux_signals[0][2][22] , 
        \s_mux_signals[0][2][21] , \s_mux_signals[0][2][20] , 
        \s_mux_signals[0][2][19] , \s_mux_signals[0][2][18] , 
        \s_mux_signals[0][2][17] , \s_mux_signals[0][2][16] , 
        \s_mux_signals[0][2][15] , \s_mux_signals[0][2][14] , 
        \s_mux_signals[0][2][13] , \s_mux_signals[0][2][12] , 
        \s_mux_signals[0][2][11] , \s_mux_signals[0][2][10] , 
        \s_mux_signals[0][2][9] , \s_mux_signals[0][2][8] , 
        \s_mux_signals[0][2][7] , \s_mux_signals[0][2][6] , 
        \s_mux_signals[0][2][5] , \s_mux_signals[0][2][4] , 
        \s_mux_signals[0][2][3] , \s_mux_signals[0][2][2] , 
        \s_mux_signals[0][2][1] , \s_mux_signals[0][2][0] }) );
  NRegister_N32_72 TargReg_i_3 ( .clk(BTB_clk), .reset(n330), .data_in({n124, 
        n120, n117, n114, n111, n108, n105, n102, n99, n96, n93, n90, n87, n84, 
        n81, n78, n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, 
        n39, n36, n33, n30}), .enable(n19), .load(s_regenabl_target[28]), 
        .data_out({\s_mux_signals[0][3][31] , \s_mux_signals[0][3][30] , 
        \s_mux_signals[0][3][29] , \s_mux_signals[0][3][28] , 
        \s_mux_signals[0][3][27] , \s_mux_signals[0][3][26] , 
        \s_mux_signals[0][3][25] , \s_mux_signals[0][3][24] , 
        \s_mux_signals[0][3][23] , \s_mux_signals[0][3][22] , 
        \s_mux_signals[0][3][21] , \s_mux_signals[0][3][20] , 
        \s_mux_signals[0][3][19] , \s_mux_signals[0][3][18] , 
        \s_mux_signals[0][3][17] , \s_mux_signals[0][3][16] , 
        \s_mux_signals[0][3][15] , \s_mux_signals[0][3][14] , 
        \s_mux_signals[0][3][13] , \s_mux_signals[0][3][12] , 
        \s_mux_signals[0][3][11] , \s_mux_signals[0][3][10] , 
        \s_mux_signals[0][3][9] , \s_mux_signals[0][3][8] , 
        \s_mux_signals[0][3][7] , \s_mux_signals[0][3][6] , 
        \s_mux_signals[0][3][5] , \s_mux_signals[0][3][4] , 
        \s_mux_signals[0][3][3] , \s_mux_signals[0][3][2] , 
        \s_mux_signals[0][3][1] , \s_mux_signals[0][3][0] }) );
  NRegister_N32_71 TargReg_i_4 ( .clk(BTB_clk), .reset(n330), .data_in({n124, 
        n120, n117, n114, n111, n108, n105, n102, n99, n96, n93, n90, n87, n84, 
        n81, n78, n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, 
        n39, n36, n33, n30}), .enable(n20), .load(s_regenabl_target[27]), 
        .data_out({\s_mux_signals[0][4][31] , \s_mux_signals[0][4][30] , 
        \s_mux_signals[0][4][29] , \s_mux_signals[0][4][28] , 
        \s_mux_signals[0][4][27] , \s_mux_signals[0][4][26] , 
        \s_mux_signals[0][4][25] , \s_mux_signals[0][4][24] , 
        \s_mux_signals[0][4][23] , \s_mux_signals[0][4][22] , 
        \s_mux_signals[0][4][21] , \s_mux_signals[0][4][20] , 
        \s_mux_signals[0][4][19] , \s_mux_signals[0][4][18] , 
        \s_mux_signals[0][4][17] , \s_mux_signals[0][4][16] , 
        \s_mux_signals[0][4][15] , \s_mux_signals[0][4][14] , 
        \s_mux_signals[0][4][13] , \s_mux_signals[0][4][12] , 
        \s_mux_signals[0][4][11] , \s_mux_signals[0][4][10] , 
        \s_mux_signals[0][4][9] , \s_mux_signals[0][4][8] , 
        \s_mux_signals[0][4][7] , \s_mux_signals[0][4][6] , 
        \s_mux_signals[0][4][5] , \s_mux_signals[0][4][4] , 
        \s_mux_signals[0][4][3] , \s_mux_signals[0][4][2] , 
        \s_mux_signals[0][4][1] , \s_mux_signals[0][4][0] }) );
  NRegister_N32_70 TargReg_i_5 ( .clk(BTB_clk), .reset(n330), .data_in({n124, 
        n120, n117, n114, n111, n108, n105, n102, n99, n96, n93, n90, n87, n84, 
        n81, n78, n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, 
        n39, n36, n33, n30}), .enable(n20), .load(s_regenabl_target[26]), 
        .data_out({\s_mux_signals[0][5][31] , \s_mux_signals[0][5][30] , 
        \s_mux_signals[0][5][29] , \s_mux_signals[0][5][28] , 
        \s_mux_signals[0][5][27] , \s_mux_signals[0][5][26] , 
        \s_mux_signals[0][5][25] , \s_mux_signals[0][5][24] , 
        \s_mux_signals[0][5][23] , \s_mux_signals[0][5][22] , 
        \s_mux_signals[0][5][21] , \s_mux_signals[0][5][20] , 
        \s_mux_signals[0][5][19] , \s_mux_signals[0][5][18] , 
        \s_mux_signals[0][5][17] , \s_mux_signals[0][5][16] , 
        \s_mux_signals[0][5][15] , \s_mux_signals[0][5][14] , 
        \s_mux_signals[0][5][13] , \s_mux_signals[0][5][12] , 
        \s_mux_signals[0][5][11] , \s_mux_signals[0][5][10] , 
        \s_mux_signals[0][5][9] , \s_mux_signals[0][5][8] , 
        \s_mux_signals[0][5][7] , \s_mux_signals[0][5][6] , 
        \s_mux_signals[0][5][5] , \s_mux_signals[0][5][4] , 
        \s_mux_signals[0][5][3] , \s_mux_signals[0][5][2] , 
        \s_mux_signals[0][5][1] , \s_mux_signals[0][5][0] }) );
  NRegister_N32_69 TargReg_i_6 ( .clk(BTB_clk), .reset(n330), .data_in({n125, 
        n120, n117, n114, n111, n108, n105, n102, n99, n96, n93, n90, n87, n84, 
        n81, n78, n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, 
        n39, n36, n33, n30}), .enable(n20), .load(s_regenabl_target[25]), 
        .data_out({\s_mux_signals[0][6][31] , \s_mux_signals[0][6][30] , 
        \s_mux_signals[0][6][29] , \s_mux_signals[0][6][28] , 
        \s_mux_signals[0][6][27] , \s_mux_signals[0][6][26] , 
        \s_mux_signals[0][6][25] , \s_mux_signals[0][6][24] , 
        \s_mux_signals[0][6][23] , \s_mux_signals[0][6][22] , 
        \s_mux_signals[0][6][21] , \s_mux_signals[0][6][20] , 
        \s_mux_signals[0][6][19] , \s_mux_signals[0][6][18] , 
        \s_mux_signals[0][6][17] , \s_mux_signals[0][6][16] , 
        \s_mux_signals[0][6][15] , \s_mux_signals[0][6][14] , 
        \s_mux_signals[0][6][13] , \s_mux_signals[0][6][12] , 
        \s_mux_signals[0][6][11] , \s_mux_signals[0][6][10] , 
        \s_mux_signals[0][6][9] , \s_mux_signals[0][6][8] , 
        \s_mux_signals[0][6][7] , \s_mux_signals[0][6][6] , 
        \s_mux_signals[0][6][5] , \s_mux_signals[0][6][4] , 
        \s_mux_signals[0][6][3] , \s_mux_signals[0][6][2] , 
        \s_mux_signals[0][6][1] , \s_mux_signals[0][6][0] }) );
  NRegister_N32_68 TargReg_i_7 ( .clk(BTB_clk), .reset(n330), .data_in({n124, 
        n120, n117, n114, n111, n108, n105, n102, n99, n96, n93, n90, n87, n84, 
        n81, n78, n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, 
        n39, n36, n33, n30}), .enable(n20), .load(s_regenabl_target[24]), 
        .data_out({\s_mux_signals[0][7][31] , \s_mux_signals[0][7][30] , 
        \s_mux_signals[0][7][29] , \s_mux_signals[0][7][28] , 
        \s_mux_signals[0][7][27] , \s_mux_signals[0][7][26] , 
        \s_mux_signals[0][7][25] , \s_mux_signals[0][7][24] , 
        \s_mux_signals[0][7][23] , \s_mux_signals[0][7][22] , 
        \s_mux_signals[0][7][21] , \s_mux_signals[0][7][20] , 
        \s_mux_signals[0][7][19] , \s_mux_signals[0][7][18] , 
        \s_mux_signals[0][7][17] , \s_mux_signals[0][7][16] , 
        \s_mux_signals[0][7][15] , \s_mux_signals[0][7][14] , 
        \s_mux_signals[0][7][13] , \s_mux_signals[0][7][12] , 
        \s_mux_signals[0][7][11] , \s_mux_signals[0][7][10] , 
        \s_mux_signals[0][7][9] , \s_mux_signals[0][7][8] , 
        \s_mux_signals[0][7][7] , \s_mux_signals[0][7][6] , 
        \s_mux_signals[0][7][5] , \s_mux_signals[0][7][4] , 
        \s_mux_signals[0][7][3] , \s_mux_signals[0][7][2] , 
        \s_mux_signals[0][7][1] , \s_mux_signals[0][7][0] }) );
  NRegister_N32_67 TargReg_i_8 ( .clk(BTB_clk), .reset(n330), .data_in({n125, 
        n120, n117, n114, n111, n108, n105, n102, n99, n96, n93, n90, n87, n84, 
        n81, n78, n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, 
        n39, n36, n33, n30}), .enable(n20), .load(s_regenabl_target[23]), 
        .data_out({\s_mux_signals[0][8][31] , \s_mux_signals[0][8][30] , 
        \s_mux_signals[0][8][29] , \s_mux_signals[0][8][28] , 
        \s_mux_signals[0][8][27] , \s_mux_signals[0][8][26] , 
        \s_mux_signals[0][8][25] , \s_mux_signals[0][8][24] , 
        \s_mux_signals[0][8][23] , \s_mux_signals[0][8][22] , 
        \s_mux_signals[0][8][21] , \s_mux_signals[0][8][20] , 
        \s_mux_signals[0][8][19] , \s_mux_signals[0][8][18] , 
        \s_mux_signals[0][8][17] , \s_mux_signals[0][8][16] , 
        \s_mux_signals[0][8][15] , \s_mux_signals[0][8][14] , 
        \s_mux_signals[0][8][13] , \s_mux_signals[0][8][12] , 
        \s_mux_signals[0][8][11] , \s_mux_signals[0][8][10] , 
        \s_mux_signals[0][8][9] , \s_mux_signals[0][8][8] , 
        \s_mux_signals[0][8][7] , \s_mux_signals[0][8][6] , 
        \s_mux_signals[0][8][5] , \s_mux_signals[0][8][4] , 
        \s_mux_signals[0][8][3] , \s_mux_signals[0][8][2] , 
        \s_mux_signals[0][8][1] , \s_mux_signals[0][8][0] }) );
  NRegister_N32_66 TargReg_i_9 ( .clk(BTB_clk), .reset(n329), .data_in({n124, 
        n120, n117, n114, n111, n108, n105, n102, n99, n96, n93, n90, n87, n84, 
        n81, n78, n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, 
        n39, n36, n33, n30}), .enable(n20), .load(s_regenabl_target[22]), 
        .data_out({\s_mux_signals[0][9][31] , \s_mux_signals[0][9][30] , 
        \s_mux_signals[0][9][29] , \s_mux_signals[0][9][28] , 
        \s_mux_signals[0][9][27] , \s_mux_signals[0][9][26] , 
        \s_mux_signals[0][9][25] , \s_mux_signals[0][9][24] , 
        \s_mux_signals[0][9][23] , \s_mux_signals[0][9][22] , 
        \s_mux_signals[0][9][21] , \s_mux_signals[0][9][20] , 
        \s_mux_signals[0][9][19] , \s_mux_signals[0][9][18] , 
        \s_mux_signals[0][9][17] , \s_mux_signals[0][9][16] , 
        \s_mux_signals[0][9][15] , \s_mux_signals[0][9][14] , 
        \s_mux_signals[0][9][13] , \s_mux_signals[0][9][12] , 
        \s_mux_signals[0][9][11] , \s_mux_signals[0][9][10] , 
        \s_mux_signals[0][9][9] , \s_mux_signals[0][9][8] , 
        \s_mux_signals[0][9][7] , \s_mux_signals[0][9][6] , 
        \s_mux_signals[0][9][5] , \s_mux_signals[0][9][4] , 
        \s_mux_signals[0][9][3] , \s_mux_signals[0][9][2] , 
        \s_mux_signals[0][9][1] , \s_mux_signals[0][9][0] }) );
  NRegister_N32_65 TargReg_i_10 ( .clk(BTB_clk), .reset(n329), .data_in({n124, 
        n120, n117, n114, n111, n108, n105, n102, n99, n96, n93, n90, n87, n84, 
        n81, n78, n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, 
        n39, n36, n33, n30}), .enable(n20), .load(s_regenabl_target[21]), 
        .data_out({\s_mux_signals[0][10][31] , \s_mux_signals[0][10][30] , 
        \s_mux_signals[0][10][29] , \s_mux_signals[0][10][28] , 
        \s_mux_signals[0][10][27] , \s_mux_signals[0][10][26] , 
        \s_mux_signals[0][10][25] , \s_mux_signals[0][10][24] , 
        \s_mux_signals[0][10][23] , \s_mux_signals[0][10][22] , 
        \s_mux_signals[0][10][21] , \s_mux_signals[0][10][20] , 
        \s_mux_signals[0][10][19] , \s_mux_signals[0][10][18] , 
        \s_mux_signals[0][10][17] , \s_mux_signals[0][10][16] , 
        \s_mux_signals[0][10][15] , \s_mux_signals[0][10][14] , 
        \s_mux_signals[0][10][13] , \s_mux_signals[0][10][12] , 
        \s_mux_signals[0][10][11] , \s_mux_signals[0][10][10] , 
        \s_mux_signals[0][10][9] , \s_mux_signals[0][10][8] , 
        \s_mux_signals[0][10][7] , \s_mux_signals[0][10][6] , 
        \s_mux_signals[0][10][5] , \s_mux_signals[0][10][4] , 
        \s_mux_signals[0][10][3] , \s_mux_signals[0][10][2] , 
        \s_mux_signals[0][10][1] , \s_mux_signals[0][10][0] }) );
  NRegister_N32_64 TargReg_i_11 ( .clk(BTB_clk), .reset(n329), .data_in({n125, 
        n120, n117, n114, n111, n108, n105, n102, n99, n96, n93, n90, n87, n84, 
        n81, n78, n75, n72, n69, n66, n63, n60, n57, n54, n51, n48, n45, n42, 
        n39, n36, n33, n30}), .enable(n20), .load(s_regenabl_target[20]), 
        .data_out({\s_mux_signals[0][11][31] , \s_mux_signals[0][11][30] , 
        \s_mux_signals[0][11][29] , \s_mux_signals[0][11][28] , 
        \s_mux_signals[0][11][27] , \s_mux_signals[0][11][26] , 
        \s_mux_signals[0][11][25] , \s_mux_signals[0][11][24] , 
        \s_mux_signals[0][11][23] , \s_mux_signals[0][11][22] , 
        \s_mux_signals[0][11][21] , \s_mux_signals[0][11][20] , 
        \s_mux_signals[0][11][19] , \s_mux_signals[0][11][18] , 
        \s_mux_signals[0][11][17] , \s_mux_signals[0][11][16] , 
        \s_mux_signals[0][11][15] , \s_mux_signals[0][11][14] , 
        \s_mux_signals[0][11][13] , \s_mux_signals[0][11][12] , 
        \s_mux_signals[0][11][11] , \s_mux_signals[0][11][10] , 
        \s_mux_signals[0][11][9] , \s_mux_signals[0][11][8] , 
        \s_mux_signals[0][11][7] , \s_mux_signals[0][11][6] , 
        \s_mux_signals[0][11][5] , \s_mux_signals[0][11][4] , 
        \s_mux_signals[0][11][3] , \s_mux_signals[0][11][2] , 
        \s_mux_signals[0][11][1] , \s_mux_signals[0][11][0] }) );
  NRegister_N32_63 TargReg_i_12 ( .clk(BTB_clk), .reset(n329), .data_in({n123, 
        n121, n118, n115, n112, n109, n106, n103, n100, n97, n94, n91, n88, 
        n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, n46, 
        n43, n40, n37, n34, n31}), .enable(n20), .load(s_regenabl_target[19]), 
        .data_out({\s_mux_signals[0][12][31] , \s_mux_signals[0][12][30] , 
        \s_mux_signals[0][12][29] , \s_mux_signals[0][12][28] , 
        \s_mux_signals[0][12][27] , \s_mux_signals[0][12][26] , 
        \s_mux_signals[0][12][25] , \s_mux_signals[0][12][24] , 
        \s_mux_signals[0][12][23] , \s_mux_signals[0][12][22] , 
        \s_mux_signals[0][12][21] , \s_mux_signals[0][12][20] , 
        \s_mux_signals[0][12][19] , \s_mux_signals[0][12][18] , 
        \s_mux_signals[0][12][17] , \s_mux_signals[0][12][16] , 
        \s_mux_signals[0][12][15] , \s_mux_signals[0][12][14] , 
        \s_mux_signals[0][12][13] , \s_mux_signals[0][12][12] , 
        \s_mux_signals[0][12][11] , \s_mux_signals[0][12][10] , 
        \s_mux_signals[0][12][9] , \s_mux_signals[0][12][8] , 
        \s_mux_signals[0][12][7] , \s_mux_signals[0][12][6] , 
        \s_mux_signals[0][12][5] , \s_mux_signals[0][12][4] , 
        \s_mux_signals[0][12][3] , \s_mux_signals[0][12][2] , 
        \s_mux_signals[0][12][1] , \s_mux_signals[0][12][0] }) );
  NRegister_N32_62 TargReg_i_13 ( .clk(BTB_clk), .reset(n329), .data_in({n123, 
        n121, n118, n115, n112, n109, n106, n103, n100, n97, n94, n91, n88, 
        n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, n46, 
        n43, n40, n37, n34, n31}), .enable(n20), .load(s_regenabl_target[18]), 
        .data_out({\s_mux_signals[0][13][31] , \s_mux_signals[0][13][30] , 
        \s_mux_signals[0][13][29] , \s_mux_signals[0][13][28] , 
        \s_mux_signals[0][13][27] , \s_mux_signals[0][13][26] , 
        \s_mux_signals[0][13][25] , \s_mux_signals[0][13][24] , 
        \s_mux_signals[0][13][23] , \s_mux_signals[0][13][22] , 
        \s_mux_signals[0][13][21] , \s_mux_signals[0][13][20] , 
        \s_mux_signals[0][13][19] , \s_mux_signals[0][13][18] , 
        \s_mux_signals[0][13][17] , \s_mux_signals[0][13][16] , 
        \s_mux_signals[0][13][15] , \s_mux_signals[0][13][14] , 
        \s_mux_signals[0][13][13] , \s_mux_signals[0][13][12] , 
        \s_mux_signals[0][13][11] , \s_mux_signals[0][13][10] , 
        \s_mux_signals[0][13][9] , \s_mux_signals[0][13][8] , 
        \s_mux_signals[0][13][7] , \s_mux_signals[0][13][6] , 
        \s_mux_signals[0][13][5] , \s_mux_signals[0][13][4] , 
        \s_mux_signals[0][13][3] , \s_mux_signals[0][13][2] , 
        \s_mux_signals[0][13][1] , \s_mux_signals[0][13][0] }) );
  NRegister_N32_61 TargReg_i_14 ( .clk(BTB_clk), .reset(n329), .data_in({n123, 
        n121, n118, n115, n112, n109, n106, n103, n100, n97, n94, n91, n88, 
        n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, n46, 
        n43, n40, n37, n34, n31}), .enable(n20), .load(s_regenabl_target[17]), 
        .data_out({\s_mux_signals[0][14][31] , \s_mux_signals[0][14][30] , 
        \s_mux_signals[0][14][29] , \s_mux_signals[0][14][28] , 
        \s_mux_signals[0][14][27] , \s_mux_signals[0][14][26] , 
        \s_mux_signals[0][14][25] , \s_mux_signals[0][14][24] , 
        \s_mux_signals[0][14][23] , \s_mux_signals[0][14][22] , 
        \s_mux_signals[0][14][21] , \s_mux_signals[0][14][20] , 
        \s_mux_signals[0][14][19] , \s_mux_signals[0][14][18] , 
        \s_mux_signals[0][14][17] , \s_mux_signals[0][14][16] , 
        \s_mux_signals[0][14][15] , \s_mux_signals[0][14][14] , 
        \s_mux_signals[0][14][13] , \s_mux_signals[0][14][12] , 
        \s_mux_signals[0][14][11] , \s_mux_signals[0][14][10] , 
        \s_mux_signals[0][14][9] , \s_mux_signals[0][14][8] , 
        \s_mux_signals[0][14][7] , \s_mux_signals[0][14][6] , 
        \s_mux_signals[0][14][5] , \s_mux_signals[0][14][4] , 
        \s_mux_signals[0][14][3] , \s_mux_signals[0][14][2] , 
        \s_mux_signals[0][14][1] , \s_mux_signals[0][14][0] }) );
  NRegister_N32_60 TargReg_i_15 ( .clk(BTB_clk), .reset(n329), .data_in({n123, 
        n121, n118, n115, n112, n109, n106, n103, n100, n97, n94, n91, n88, 
        n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, n46, 
        n43, n40, n37, n34, n31}), .enable(n20), .load(s_regenabl_target[16]), 
        .data_out({\s_mux_signals[0][15][31] , \s_mux_signals[0][15][30] , 
        \s_mux_signals[0][15][29] , \s_mux_signals[0][15][28] , 
        \s_mux_signals[0][15][27] , \s_mux_signals[0][15][26] , 
        \s_mux_signals[0][15][25] , \s_mux_signals[0][15][24] , 
        \s_mux_signals[0][15][23] , \s_mux_signals[0][15][22] , 
        \s_mux_signals[0][15][21] , \s_mux_signals[0][15][20] , 
        \s_mux_signals[0][15][19] , \s_mux_signals[0][15][18] , 
        \s_mux_signals[0][15][17] , \s_mux_signals[0][15][16] , 
        \s_mux_signals[0][15][15] , \s_mux_signals[0][15][14] , 
        \s_mux_signals[0][15][13] , \s_mux_signals[0][15][12] , 
        \s_mux_signals[0][15][11] , \s_mux_signals[0][15][10] , 
        \s_mux_signals[0][15][9] , \s_mux_signals[0][15][8] , 
        \s_mux_signals[0][15][7] , \s_mux_signals[0][15][6] , 
        \s_mux_signals[0][15][5] , \s_mux_signals[0][15][4] , 
        \s_mux_signals[0][15][3] , \s_mux_signals[0][15][2] , 
        \s_mux_signals[0][15][1] , \s_mux_signals[0][15][0] }) );
  NRegister_N32_59 TargReg_i_16 ( .clk(BTB_clk), .reset(n329), .data_in({n123, 
        n121, n118, n115, n112, n109, n106, n103, n100, n97, n94, n91, n88, 
        n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, n46, 
        n43, n40, n37, n34, n31}), .enable(n21), .load(s_regenabl_target[15]), 
        .data_out({\s_mux_signals[0][16][31] , \s_mux_signals[0][16][30] , 
        \s_mux_signals[0][16][29] , \s_mux_signals[0][16][28] , 
        \s_mux_signals[0][16][27] , \s_mux_signals[0][16][26] , 
        \s_mux_signals[0][16][25] , \s_mux_signals[0][16][24] , 
        \s_mux_signals[0][16][23] , \s_mux_signals[0][16][22] , 
        \s_mux_signals[0][16][21] , \s_mux_signals[0][16][20] , 
        \s_mux_signals[0][16][19] , \s_mux_signals[0][16][18] , 
        \s_mux_signals[0][16][17] , \s_mux_signals[0][16][16] , 
        \s_mux_signals[0][16][15] , \s_mux_signals[0][16][14] , 
        \s_mux_signals[0][16][13] , \s_mux_signals[0][16][12] , 
        \s_mux_signals[0][16][11] , \s_mux_signals[0][16][10] , 
        \s_mux_signals[0][16][9] , \s_mux_signals[0][16][8] , 
        \s_mux_signals[0][16][7] , \s_mux_signals[0][16][6] , 
        \s_mux_signals[0][16][5] , \s_mux_signals[0][16][4] , 
        \s_mux_signals[0][16][3] , \s_mux_signals[0][16][2] , 
        \s_mux_signals[0][16][1] , \s_mux_signals[0][16][0] }) );
  NRegister_N32_58 TargReg_i_17 ( .clk(BTB_clk), .reset(n329), .data_in({n123, 
        n121, n118, n115, n112, n109, n106, n103, n100, n97, n94, n91, n88, 
        n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, n46, 
        n43, n40, n37, n34, n31}), .enable(n21), .load(s_regenabl_target[14]), 
        .data_out({\s_mux_signals[0][17][31] , \s_mux_signals[0][17][30] , 
        \s_mux_signals[0][17][29] , \s_mux_signals[0][17][28] , 
        \s_mux_signals[0][17][27] , \s_mux_signals[0][17][26] , 
        \s_mux_signals[0][17][25] , \s_mux_signals[0][17][24] , 
        \s_mux_signals[0][17][23] , \s_mux_signals[0][17][22] , 
        \s_mux_signals[0][17][21] , \s_mux_signals[0][17][20] , 
        \s_mux_signals[0][17][19] , \s_mux_signals[0][17][18] , 
        \s_mux_signals[0][17][17] , \s_mux_signals[0][17][16] , 
        \s_mux_signals[0][17][15] , \s_mux_signals[0][17][14] , 
        \s_mux_signals[0][17][13] , \s_mux_signals[0][17][12] , 
        \s_mux_signals[0][17][11] , \s_mux_signals[0][17][10] , 
        \s_mux_signals[0][17][9] , \s_mux_signals[0][17][8] , 
        \s_mux_signals[0][17][7] , \s_mux_signals[0][17][6] , 
        \s_mux_signals[0][17][5] , \s_mux_signals[0][17][4] , 
        \s_mux_signals[0][17][3] , \s_mux_signals[0][17][2] , 
        \s_mux_signals[0][17][1] , \s_mux_signals[0][17][0] }) );
  NRegister_N32_57 TargReg_i_18 ( .clk(BTB_clk), .reset(n329), .data_in({n123, 
        n121, n118, n115, n112, n109, n106, n103, n100, n97, n94, n91, n88, 
        n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, n46, 
        n43, n40, n37, n34, n31}), .enable(n21), .load(s_regenabl_target[13]), 
        .data_out({\s_mux_signals[0][18][31] , \s_mux_signals[0][18][30] , 
        \s_mux_signals[0][18][29] , \s_mux_signals[0][18][28] , 
        \s_mux_signals[0][18][27] , \s_mux_signals[0][18][26] , 
        \s_mux_signals[0][18][25] , \s_mux_signals[0][18][24] , 
        \s_mux_signals[0][18][23] , \s_mux_signals[0][18][22] , 
        \s_mux_signals[0][18][21] , \s_mux_signals[0][18][20] , 
        \s_mux_signals[0][18][19] , \s_mux_signals[0][18][18] , 
        \s_mux_signals[0][18][17] , \s_mux_signals[0][18][16] , 
        \s_mux_signals[0][18][15] , \s_mux_signals[0][18][14] , 
        \s_mux_signals[0][18][13] , \s_mux_signals[0][18][12] , 
        \s_mux_signals[0][18][11] , \s_mux_signals[0][18][10] , 
        \s_mux_signals[0][18][9] , \s_mux_signals[0][18][8] , 
        \s_mux_signals[0][18][7] , \s_mux_signals[0][18][6] , 
        \s_mux_signals[0][18][5] , \s_mux_signals[0][18][4] , 
        \s_mux_signals[0][18][3] , \s_mux_signals[0][18][2] , 
        \s_mux_signals[0][18][1] , \s_mux_signals[0][18][0] }) );
  NRegister_N32_56 TargReg_i_19 ( .clk(BTB_clk), .reset(n329), .data_in({n123, 
        n121, n118, n115, n112, n109, n106, n103, n100, n97, n94, n91, n88, 
        n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, n46, 
        n43, n40, n37, n34, n31}), .enable(n21), .load(s_regenabl_target[12]), 
        .data_out({\s_mux_signals[0][19][31] , \s_mux_signals[0][19][30] , 
        \s_mux_signals[0][19][29] , \s_mux_signals[0][19][28] , 
        \s_mux_signals[0][19][27] , \s_mux_signals[0][19][26] , 
        \s_mux_signals[0][19][25] , \s_mux_signals[0][19][24] , 
        \s_mux_signals[0][19][23] , \s_mux_signals[0][19][22] , 
        \s_mux_signals[0][19][21] , \s_mux_signals[0][19][20] , 
        \s_mux_signals[0][19][19] , \s_mux_signals[0][19][18] , 
        \s_mux_signals[0][19][17] , \s_mux_signals[0][19][16] , 
        \s_mux_signals[0][19][15] , \s_mux_signals[0][19][14] , 
        \s_mux_signals[0][19][13] , \s_mux_signals[0][19][12] , 
        \s_mux_signals[0][19][11] , \s_mux_signals[0][19][10] , 
        \s_mux_signals[0][19][9] , \s_mux_signals[0][19][8] , 
        \s_mux_signals[0][19][7] , \s_mux_signals[0][19][6] , 
        \s_mux_signals[0][19][5] , \s_mux_signals[0][19][4] , 
        \s_mux_signals[0][19][3] , \s_mux_signals[0][19][2] , 
        \s_mux_signals[0][19][1] , \s_mux_signals[0][19][0] }) );
  NRegister_N32_55 TargReg_i_20 ( .clk(BTB_clk), .reset(n329), .data_in({n123, 
        n121, n118, n115, n112, n109, n106, n103, n100, n97, n94, n91, n88, 
        n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, n46, 
        n43, n40, n37, n34, n31}), .enable(n21), .load(s_regenabl_target[11]), 
        .data_out({\s_mux_signals[0][20][31] , \s_mux_signals[0][20][30] , 
        \s_mux_signals[0][20][29] , \s_mux_signals[0][20][28] , 
        \s_mux_signals[0][20][27] , \s_mux_signals[0][20][26] , 
        \s_mux_signals[0][20][25] , \s_mux_signals[0][20][24] , 
        \s_mux_signals[0][20][23] , \s_mux_signals[0][20][22] , 
        \s_mux_signals[0][20][21] , \s_mux_signals[0][20][20] , 
        \s_mux_signals[0][20][19] , \s_mux_signals[0][20][18] , 
        \s_mux_signals[0][20][17] , \s_mux_signals[0][20][16] , 
        \s_mux_signals[0][20][15] , \s_mux_signals[0][20][14] , 
        \s_mux_signals[0][20][13] , \s_mux_signals[0][20][12] , 
        \s_mux_signals[0][20][11] , \s_mux_signals[0][20][10] , 
        \s_mux_signals[0][20][9] , \s_mux_signals[0][20][8] , 
        \s_mux_signals[0][20][7] , \s_mux_signals[0][20][6] , 
        \s_mux_signals[0][20][5] , \s_mux_signals[0][20][4] , 
        \s_mux_signals[0][20][3] , \s_mux_signals[0][20][2] , 
        \s_mux_signals[0][20][1] , \s_mux_signals[0][20][0] }) );
  NRegister_N32_54 TargReg_i_21 ( .clk(BTB_clk), .reset(n328), .data_in({n123, 
        n121, n118, n115, n112, n109, n106, n103, n100, n97, n94, n91, n88, 
        n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, n46, 
        n43, n40, n37, n34, n31}), .enable(n21), .load(s_regenabl_target[10]), 
        .data_out({\s_mux_signals[0][21][31] , \s_mux_signals[0][21][30] , 
        \s_mux_signals[0][21][29] , \s_mux_signals[0][21][28] , 
        \s_mux_signals[0][21][27] , \s_mux_signals[0][21][26] , 
        \s_mux_signals[0][21][25] , \s_mux_signals[0][21][24] , 
        \s_mux_signals[0][21][23] , \s_mux_signals[0][21][22] , 
        \s_mux_signals[0][21][21] , \s_mux_signals[0][21][20] , 
        \s_mux_signals[0][21][19] , \s_mux_signals[0][21][18] , 
        \s_mux_signals[0][21][17] , \s_mux_signals[0][21][16] , 
        \s_mux_signals[0][21][15] , \s_mux_signals[0][21][14] , 
        \s_mux_signals[0][21][13] , \s_mux_signals[0][21][12] , 
        \s_mux_signals[0][21][11] , \s_mux_signals[0][21][10] , 
        \s_mux_signals[0][21][9] , \s_mux_signals[0][21][8] , 
        \s_mux_signals[0][21][7] , \s_mux_signals[0][21][6] , 
        \s_mux_signals[0][21][5] , \s_mux_signals[0][21][4] , 
        \s_mux_signals[0][21][3] , \s_mux_signals[0][21][2] , 
        \s_mux_signals[0][21][1] , \s_mux_signals[0][21][0] }) );
  NRegister_N32_53 TargReg_i_22 ( .clk(BTB_clk), .reset(n328), .data_in({n125, 
        n121, n118, n115, n112, n109, n106, n103, n100, n97, n94, n91, n88, 
        n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, n46, 
        n43, n40, n37, n34, n31}), .enable(n21), .load(s_regenabl_target[9]), 
        .data_out({\s_mux_signals[0][22][31] , \s_mux_signals[0][22][30] , 
        \s_mux_signals[0][22][29] , \s_mux_signals[0][22][28] , 
        \s_mux_signals[0][22][27] , \s_mux_signals[0][22][26] , 
        \s_mux_signals[0][22][25] , \s_mux_signals[0][22][24] , 
        \s_mux_signals[0][22][23] , \s_mux_signals[0][22][22] , 
        \s_mux_signals[0][22][21] , \s_mux_signals[0][22][20] , 
        \s_mux_signals[0][22][19] , \s_mux_signals[0][22][18] , 
        \s_mux_signals[0][22][17] , \s_mux_signals[0][22][16] , 
        \s_mux_signals[0][22][15] , \s_mux_signals[0][22][14] , 
        \s_mux_signals[0][22][13] , \s_mux_signals[0][22][12] , 
        \s_mux_signals[0][22][11] , \s_mux_signals[0][22][10] , 
        \s_mux_signals[0][22][9] , \s_mux_signals[0][22][8] , 
        \s_mux_signals[0][22][7] , \s_mux_signals[0][22][6] , 
        \s_mux_signals[0][22][5] , \s_mux_signals[0][22][4] , 
        \s_mux_signals[0][22][3] , \s_mux_signals[0][22][2] , 
        \s_mux_signals[0][22][1] , \s_mux_signals[0][22][0] }) );
  NRegister_N32_52 TargReg_i_23 ( .clk(BTB_clk), .reset(n328), .data_in({n123, 
        n121, n118, n115, n112, n109, n106, n103, n100, n97, n94, n91, n88, 
        n85, n82, n79, n76, n73, n70, n67, n64, n61, n58, n55, n52, n49, n46, 
        n43, n40, n37, n34, n31}), .enable(n21), .load(s_regenabl_target[8]), 
        .data_out({\s_mux_signals[0][23][31] , \s_mux_signals[0][23][30] , 
        \s_mux_signals[0][23][29] , \s_mux_signals[0][23][28] , 
        \s_mux_signals[0][23][27] , \s_mux_signals[0][23][26] , 
        \s_mux_signals[0][23][25] , \s_mux_signals[0][23][24] , 
        \s_mux_signals[0][23][23] , \s_mux_signals[0][23][22] , 
        \s_mux_signals[0][23][21] , \s_mux_signals[0][23][20] , 
        \s_mux_signals[0][23][19] , \s_mux_signals[0][23][18] , 
        \s_mux_signals[0][23][17] , \s_mux_signals[0][23][16] , 
        \s_mux_signals[0][23][15] , \s_mux_signals[0][23][14] , 
        \s_mux_signals[0][23][13] , \s_mux_signals[0][23][12] , 
        \s_mux_signals[0][23][11] , \s_mux_signals[0][23][10] , 
        \s_mux_signals[0][23][9] , \s_mux_signals[0][23][8] , 
        \s_mux_signals[0][23][7] , \s_mux_signals[0][23][6] , 
        \s_mux_signals[0][23][5] , \s_mux_signals[0][23][4] , 
        \s_mux_signals[0][23][3] , \s_mux_signals[0][23][2] , 
        \s_mux_signals[0][23][1] , \s_mux_signals[0][23][0] }) );
  NRegister_N32_51 TargReg_i_24 ( .clk(BTB_clk), .reset(n328), .data_in({n124, 
        n122, n119, n116, n113, n110, n107, n104, n101, n98, n95, n92, n89, 
        n86, n83, n80, n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, 
        n44, n41, n38, n35, n32}), .enable(n21), .load(s_regenabl_target[7]), 
        .data_out({\s_mux_signals[0][24][31] , \s_mux_signals[0][24][30] , 
        \s_mux_signals[0][24][29] , \s_mux_signals[0][24][28] , 
        \s_mux_signals[0][24][27] , \s_mux_signals[0][24][26] , 
        \s_mux_signals[0][24][25] , \s_mux_signals[0][24][24] , 
        \s_mux_signals[0][24][23] , \s_mux_signals[0][24][22] , 
        \s_mux_signals[0][24][21] , \s_mux_signals[0][24][20] , 
        \s_mux_signals[0][24][19] , \s_mux_signals[0][24][18] , 
        \s_mux_signals[0][24][17] , \s_mux_signals[0][24][16] , 
        \s_mux_signals[0][24][15] , \s_mux_signals[0][24][14] , 
        \s_mux_signals[0][24][13] , \s_mux_signals[0][24][12] , 
        \s_mux_signals[0][24][11] , \s_mux_signals[0][24][10] , 
        \s_mux_signals[0][24][9] , \s_mux_signals[0][24][8] , 
        \s_mux_signals[0][24][7] , \s_mux_signals[0][24][6] , 
        \s_mux_signals[0][24][5] , \s_mux_signals[0][24][4] , 
        \s_mux_signals[0][24][3] , \s_mux_signals[0][24][2] , 
        \s_mux_signals[0][24][1] , \s_mux_signals[0][24][0] }) );
  NRegister_N32_50 TargReg_i_25 ( .clk(BTB_clk), .reset(n328), .data_in({n124, 
        n122, n119, n116, n113, n110, n107, n104, n101, n98, n95, n92, n89, 
        n86, n83, n80, n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, 
        n44, n41, n38, n35, n32}), .enable(n21), .load(s_regenabl_target[6]), 
        .data_out({\s_mux_signals[0][25][31] , \s_mux_signals[0][25][30] , 
        \s_mux_signals[0][25][29] , \s_mux_signals[0][25][28] , 
        \s_mux_signals[0][25][27] , \s_mux_signals[0][25][26] , 
        \s_mux_signals[0][25][25] , \s_mux_signals[0][25][24] , 
        \s_mux_signals[0][25][23] , \s_mux_signals[0][25][22] , 
        \s_mux_signals[0][25][21] , \s_mux_signals[0][25][20] , 
        \s_mux_signals[0][25][19] , \s_mux_signals[0][25][18] , 
        \s_mux_signals[0][25][17] , \s_mux_signals[0][25][16] , 
        \s_mux_signals[0][25][15] , \s_mux_signals[0][25][14] , 
        \s_mux_signals[0][25][13] , \s_mux_signals[0][25][12] , 
        \s_mux_signals[0][25][11] , \s_mux_signals[0][25][10] , 
        \s_mux_signals[0][25][9] , \s_mux_signals[0][25][8] , 
        \s_mux_signals[0][25][7] , \s_mux_signals[0][25][6] , 
        \s_mux_signals[0][25][5] , \s_mux_signals[0][25][4] , 
        \s_mux_signals[0][25][3] , \s_mux_signals[0][25][2] , 
        \s_mux_signals[0][25][1] , \s_mux_signals[0][25][0] }) );
  NRegister_N32_49 TargReg_i_26 ( .clk(BTB_clk), .reset(n328), .data_in({n125, 
        n122, n119, n116, n113, n110, n107, n104, n101, n98, n95, n92, n89, 
        n86, n83, n80, n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, 
        n44, n41, n38, n35, n32}), .enable(n21), .load(s_regenabl_target[5]), 
        .data_out({\s_mux_signals[0][26][31] , \s_mux_signals[0][26][30] , 
        \s_mux_signals[0][26][29] , \s_mux_signals[0][26][28] , 
        \s_mux_signals[0][26][27] , \s_mux_signals[0][26][26] , 
        \s_mux_signals[0][26][25] , \s_mux_signals[0][26][24] , 
        \s_mux_signals[0][26][23] , \s_mux_signals[0][26][22] , 
        \s_mux_signals[0][26][21] , \s_mux_signals[0][26][20] , 
        \s_mux_signals[0][26][19] , \s_mux_signals[0][26][18] , 
        \s_mux_signals[0][26][17] , \s_mux_signals[0][26][16] , 
        \s_mux_signals[0][26][15] , \s_mux_signals[0][26][14] , 
        \s_mux_signals[0][26][13] , \s_mux_signals[0][26][12] , 
        \s_mux_signals[0][26][11] , \s_mux_signals[0][26][10] , 
        \s_mux_signals[0][26][9] , \s_mux_signals[0][26][8] , 
        \s_mux_signals[0][26][7] , \s_mux_signals[0][26][6] , 
        \s_mux_signals[0][26][5] , \s_mux_signals[0][26][4] , 
        \s_mux_signals[0][26][3] , \s_mux_signals[0][26][2] , 
        \s_mux_signals[0][26][1] , \s_mux_signals[0][26][0] }) );
  NRegister_N32_48 TargReg_i_27 ( .clk(BTB_clk), .reset(n328), .data_in({n125, 
        n122, n119, n116, n113, n110, n107, n104, n101, n98, n95, n92, n89, 
        n86, n83, n80, n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, 
        n44, n41, n38, n35, n32}), .enable(n21), .load(s_regenabl_target[4]), 
        .data_out({\s_mux_signals[0][27][31] , \s_mux_signals[0][27][30] , 
        \s_mux_signals[0][27][29] , \s_mux_signals[0][27][28] , 
        \s_mux_signals[0][27][27] , \s_mux_signals[0][27][26] , 
        \s_mux_signals[0][27][25] , \s_mux_signals[0][27][24] , 
        \s_mux_signals[0][27][23] , \s_mux_signals[0][27][22] , 
        \s_mux_signals[0][27][21] , \s_mux_signals[0][27][20] , 
        \s_mux_signals[0][27][19] , \s_mux_signals[0][27][18] , 
        \s_mux_signals[0][27][17] , \s_mux_signals[0][27][16] , 
        \s_mux_signals[0][27][15] , \s_mux_signals[0][27][14] , 
        \s_mux_signals[0][27][13] , \s_mux_signals[0][27][12] , 
        \s_mux_signals[0][27][11] , \s_mux_signals[0][27][10] , 
        \s_mux_signals[0][27][9] , \s_mux_signals[0][27][8] , 
        \s_mux_signals[0][27][7] , \s_mux_signals[0][27][6] , 
        \s_mux_signals[0][27][5] , \s_mux_signals[0][27][4] , 
        \s_mux_signals[0][27][3] , \s_mux_signals[0][27][2] , 
        \s_mux_signals[0][27][1] , \s_mux_signals[0][27][0] }) );
  NRegister_N32_47 TargReg_i_28 ( .clk(BTB_clk), .reset(n328), .data_in({n124, 
        n122, n119, n116, n113, n110, n107, n104, n101, n98, n95, n92, n89, 
        n86, n83, n80, n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, 
        n44, n41, n38, n35, n32}), .enable(n22), .load(s_regenabl_target[3]), 
        .data_out({\s_mux_signals[0][28][31] , \s_mux_signals[0][28][30] , 
        \s_mux_signals[0][28][29] , \s_mux_signals[0][28][28] , 
        \s_mux_signals[0][28][27] , \s_mux_signals[0][28][26] , 
        \s_mux_signals[0][28][25] , \s_mux_signals[0][28][24] , 
        \s_mux_signals[0][28][23] , \s_mux_signals[0][28][22] , 
        \s_mux_signals[0][28][21] , \s_mux_signals[0][28][20] , 
        \s_mux_signals[0][28][19] , \s_mux_signals[0][28][18] , 
        \s_mux_signals[0][28][17] , \s_mux_signals[0][28][16] , 
        \s_mux_signals[0][28][15] , \s_mux_signals[0][28][14] , 
        \s_mux_signals[0][28][13] , \s_mux_signals[0][28][12] , 
        \s_mux_signals[0][28][11] , \s_mux_signals[0][28][10] , 
        \s_mux_signals[0][28][9] , \s_mux_signals[0][28][8] , 
        \s_mux_signals[0][28][7] , \s_mux_signals[0][28][6] , 
        \s_mux_signals[0][28][5] , \s_mux_signals[0][28][4] , 
        \s_mux_signals[0][28][3] , \s_mux_signals[0][28][2] , 
        \s_mux_signals[0][28][1] , \s_mux_signals[0][28][0] }) );
  NRegister_N32_46 TargReg_i_29 ( .clk(BTB_clk), .reset(n328), .data_in({n125, 
        n122, n119, n116, n113, n110, n107, n104, n101, n98, n95, n92, n89, 
        n86, n83, n80, n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, 
        n44, n41, n38, n35, n32}), .enable(n22), .load(s_regenabl_target[2]), 
        .data_out({\s_mux_signals[0][29][31] , \s_mux_signals[0][29][30] , 
        \s_mux_signals[0][29][29] , \s_mux_signals[0][29][28] , 
        \s_mux_signals[0][29][27] , \s_mux_signals[0][29][26] , 
        \s_mux_signals[0][29][25] , \s_mux_signals[0][29][24] , 
        \s_mux_signals[0][29][23] , \s_mux_signals[0][29][22] , 
        \s_mux_signals[0][29][21] , \s_mux_signals[0][29][20] , 
        \s_mux_signals[0][29][19] , \s_mux_signals[0][29][18] , 
        \s_mux_signals[0][29][17] , \s_mux_signals[0][29][16] , 
        \s_mux_signals[0][29][15] , \s_mux_signals[0][29][14] , 
        \s_mux_signals[0][29][13] , \s_mux_signals[0][29][12] , 
        \s_mux_signals[0][29][11] , \s_mux_signals[0][29][10] , 
        \s_mux_signals[0][29][9] , \s_mux_signals[0][29][8] , 
        \s_mux_signals[0][29][7] , \s_mux_signals[0][29][6] , 
        \s_mux_signals[0][29][5] , \s_mux_signals[0][29][4] , 
        \s_mux_signals[0][29][3] , \s_mux_signals[0][29][2] , 
        \s_mux_signals[0][29][1] , \s_mux_signals[0][29][0] }) );
  NRegister_N32_45 TargReg_i_30 ( .clk(BTB_clk), .reset(n328), .data_in({n124, 
        n122, n119, n116, n113, n110, n107, n104, n101, n98, n95, n92, n89, 
        n86, n83, n80, n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, 
        n44, n41, n38, n35, n32}), .enable(n22), .load(s_regenabl_target[1]), 
        .data_out({\s_mux_signals[0][30][31] , \s_mux_signals[0][30][30] , 
        \s_mux_signals[0][30][29] , \s_mux_signals[0][30][28] , 
        \s_mux_signals[0][30][27] , \s_mux_signals[0][30][26] , 
        \s_mux_signals[0][30][25] , \s_mux_signals[0][30][24] , 
        \s_mux_signals[0][30][23] , \s_mux_signals[0][30][22] , 
        \s_mux_signals[0][30][21] , \s_mux_signals[0][30][20] , 
        \s_mux_signals[0][30][19] , \s_mux_signals[0][30][18] , 
        \s_mux_signals[0][30][17] , \s_mux_signals[0][30][16] , 
        \s_mux_signals[0][30][15] , \s_mux_signals[0][30][14] , 
        \s_mux_signals[0][30][13] , \s_mux_signals[0][30][12] , 
        \s_mux_signals[0][30][11] , \s_mux_signals[0][30][10] , 
        \s_mux_signals[0][30][9] , \s_mux_signals[0][30][8] , 
        \s_mux_signals[0][30][7] , \s_mux_signals[0][30][6] , 
        \s_mux_signals[0][30][5] , \s_mux_signals[0][30][4] , 
        \s_mux_signals[0][30][3] , \s_mux_signals[0][30][2] , 
        \s_mux_signals[0][30][1] , \s_mux_signals[0][30][0] }) );
  NRegister_N32_44 TargReg_i_31 ( .clk(BTB_clk), .reset(n328), .data_in({n125, 
        n122, n119, n116, n113, n110, n107, n104, n101, n98, n95, n92, n89, 
        n86, n83, n80, n77, n74, n71, n68, n65, n62, n59, n56, n53, n50, n47, 
        n44, n41, n38, n35, n32}), .enable(n22), .load(s_regenabl_target[0]), 
        .data_out({\s_mux_signals[0][31][31] , \s_mux_signals[0][31][30] , 
        \s_mux_signals[0][31][29] , \s_mux_signals[0][31][28] , 
        \s_mux_signals[0][31][27] , \s_mux_signals[0][31][26] , 
        \s_mux_signals[0][31][25] , \s_mux_signals[0][31][24] , 
        \s_mux_signals[0][31][23] , \s_mux_signals[0][31][22] , 
        \s_mux_signals[0][31][21] , \s_mux_signals[0][31][20] , 
        \s_mux_signals[0][31][19] , \s_mux_signals[0][31][18] , 
        \s_mux_signals[0][31][17] , \s_mux_signals[0][31][16] , 
        \s_mux_signals[0][31][15] , \s_mux_signals[0][31][14] , 
        \s_mux_signals[0][31][13] , \s_mux_signals[0][31][12] , 
        \s_mux_signals[0][31][11] , \s_mux_signals[0][31][10] , 
        \s_mux_signals[0][31][9] , \s_mux_signals[0][31][8] , 
        \s_mux_signals[0][31][7] , \s_mux_signals[0][31][6] , 
        \s_mux_signals[0][31][5] , \s_mux_signals[0][31][4] , 
        \s_mux_signals[0][31][3] , \s_mux_signals[0][31][2] , 
        \s_mux_signals[0][31][1] , \s_mux_signals[0][31][0] }) );
  Reg1Bit_10 HitMissReg ( .clk(BTB_clk), .reset(n335), .data_in(s_HIT_miss), 
        .enable(n320), .load(1'b1), .data_out(s_HIT_miss_Freg_Txor) );
  Reg1Bit_9 RESTORE_REG_BTB ( .clk(BTB_clk), .reset(n335), .data_in(n22), 
        .enable(n321), .load(1'b1) );
  NRotateRegister_N32 RotReg ( .clk(BTB_clk), .reset(n335), .enable(n318), 
        .load(1'b0), .data_in({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .rotate(n14), .data_out(s_regenabl_FrotateR_Tregs) );
  Mux_NBit_2x1_NBIT_IN32_124 Mux_Frot_Tentr ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .port1(s_regenabl_FrotateR_Tregs), .sel(n14), 
        .portY(s_regenabl_entry) );
  Mux_NBit_2x1_NBIT_IN32_123 Mux_Frot_Ttarg ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .port1(s_regenabl_FrotateR_Tregs), .sel(n14), 
        .portY(s_regenabl_target) );
  Mux_NBit_2x1_NBIT_IN32_122 Mux_Frot_Tsat ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .port1(s_regenabl_FrotateR_Tregs), .sel(n14), 
        .portY(s_regenabl_sat) );
  NRegister_N32_43 CompBitsReg ( .clk(BTB_clk), .reset(n328), .data_in(
        s_cmpbits_Fcmp_Tencoder), .enable(n319), .load(1'b1), .data_out(
        s_updateSat_FregCmpBits_Tsats) );
  SAT_Counter_BTB_N3_0 SAT_Cnt_i_0 ( .SAT_clk(BTB_clk), .SAT_reset(n335), 
        .SAT_enable(n318), .SAT_Ud(n28), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[0]), .SAT_setToDef(s_regenabl_sat[31]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[0]) );
  SAT_Counter_BTB_N3_31 SAT_Cnt_i_1 ( .SAT_clk(BTB_clk), .SAT_reset(n335), 
        .SAT_enable(n322), .SAT_Ud(n27), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[1]), .SAT_setToDef(s_regenabl_sat[30]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[1]) );
  SAT_Counter_BTB_N3_30 SAT_Cnt_i_2 ( .SAT_clk(BTB_clk), .SAT_reset(n335), 
        .SAT_enable(n8), .SAT_Ud(n29), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[2]), .SAT_setToDef(s_regenabl_sat[29]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[2]) );
  SAT_Counter_BTB_N3_29 SAT_Cnt_i_3 ( .SAT_clk(BTB_clk), .SAT_reset(n335), 
        .SAT_enable(n323), .SAT_Ud(n29), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[3]), .SAT_setToDef(s_regenabl_sat[28]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[3]) );
  SAT_Counter_BTB_N3_28 SAT_Cnt_i_4 ( .SAT_clk(BTB_clk), .SAT_reset(n335), 
        .SAT_enable(n318), .SAT_Ud(n29), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[4]), .SAT_setToDef(s_regenabl_sat[27]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[4]) );
  SAT_Counter_BTB_N3_27 SAT_Cnt_i_5 ( .SAT_clk(BTB_clk), .SAT_reset(n335), 
        .SAT_enable(n318), .SAT_Ud(n29), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[5]), .SAT_setToDef(s_regenabl_sat[26]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[5]) );
  SAT_Counter_BTB_N3_26 SAT_Cnt_i_6 ( .SAT_clk(BTB_clk), .SAT_reset(n335), 
        .SAT_enable(n320), .SAT_Ud(n29), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[6]), .SAT_setToDef(s_regenabl_sat[25]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[6]) );
  SAT_Counter_BTB_N3_25 SAT_Cnt_i_7 ( .SAT_clk(BTB_clk), .SAT_reset(n335), 
        .SAT_enable(n322), .SAT_Ud(n29), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[7]), .SAT_setToDef(s_regenabl_sat[24]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[7]) );
  SAT_Counter_BTB_N3_24 SAT_Cnt_i_8 ( .SAT_clk(BTB_clk), .SAT_reset(n334), 
        .SAT_enable(n321), .SAT_Ud(n29), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[8]), .SAT_setToDef(s_regenabl_sat[23]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[8]) );
  SAT_Counter_BTB_N3_23 SAT_Cnt_i_9 ( .SAT_clk(BTB_clk), .SAT_reset(n335), 
        .SAT_enable(n321), .SAT_Ud(n29), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[9]), .SAT_setToDef(s_regenabl_sat[22]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[9]) );
  SAT_Counter_BTB_N3_22 SAT_Cnt_i_10 ( .SAT_clk(BTB_clk), .SAT_reset(n335), 
        .SAT_enable(n320), .SAT_Ud(n28), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[10]), .SAT_setToDef(s_regenabl_sat[21]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[10]) );
  SAT_Counter_BTB_N3_21 SAT_Cnt_i_11 ( .SAT_clk(BTB_clk), .SAT_reset(n334), 
        .SAT_enable(n319), .SAT_Ud(n28), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[11]), .SAT_setToDef(s_regenabl_sat[20]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[11]) );
  SAT_Counter_BTB_N3_20 SAT_Cnt_i_12 ( .SAT_clk(BTB_clk), .SAT_reset(n334), 
        .SAT_enable(n322), .SAT_Ud(n28), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[12]), .SAT_setToDef(s_regenabl_sat[19]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[12]) );
  SAT_Counter_BTB_N3_19 SAT_Cnt_i_13 ( .SAT_clk(BTB_clk), .SAT_reset(n334), 
        .SAT_enable(n322), .SAT_Ud(n28), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[13]), .SAT_setToDef(s_regenabl_sat[18]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[13]) );
  SAT_Counter_BTB_N3_18 SAT_Cnt_i_14 ( .SAT_clk(BTB_clk), .SAT_reset(n334), 
        .SAT_enable(n321), .SAT_Ud(n28), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[14]), .SAT_setToDef(s_regenabl_sat[17]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[14]) );
  SAT_Counter_BTB_N3_17 SAT_Cnt_i_15 ( .SAT_clk(BTB_clk), .SAT_reset(n334), 
        .SAT_enable(n322), .SAT_Ud(n28), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[15]), .SAT_setToDef(s_regenabl_sat[16]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[15]) );
  SAT_Counter_BTB_N3_16 SAT_Cnt_i_16 ( .SAT_clk(BTB_clk), .SAT_reset(n334), 
        .SAT_enable(n319), .SAT_Ud(n28), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[16]), .SAT_setToDef(s_regenabl_sat[15]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[16]) );
  SAT_Counter_BTB_N3_15 SAT_Cnt_i_17 ( .SAT_clk(BTB_clk), .SAT_reset(n334), 
        .SAT_enable(n318), .SAT_Ud(n28), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[17]), .SAT_setToDef(s_regenabl_sat[14]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[17]) );
  SAT_Counter_BTB_N3_14 SAT_Cnt_i_18 ( .SAT_clk(BTB_clk), .SAT_reset(n333), 
        .SAT_enable(n321), .SAT_Ud(n28), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[18]), .SAT_setToDef(s_regenabl_sat[13]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[18]) );
  SAT_Counter_BTB_N3_13 SAT_Cnt_i_19 ( .SAT_clk(BTB_clk), .SAT_reset(n334), 
        .SAT_enable(n319), .SAT_Ud(n28), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[19]), .SAT_setToDef(s_regenabl_sat[12]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[19]) );
  SAT_Counter_BTB_N3_12 SAT_Cnt_i_20 ( .SAT_clk(BTB_clk), .SAT_reset(n334), 
        .SAT_enable(n8), .SAT_Ud(n28), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[20]), .SAT_setToDef(s_regenabl_sat[11]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[20]) );
  SAT_Counter_BTB_N3_11 SAT_Cnt_i_21 ( .SAT_clk(BTB_clk), .SAT_reset(n334), 
        .SAT_enable(n320), .SAT_Ud(n27), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[21]), .SAT_setToDef(s_regenabl_sat[10]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[21]) );
  SAT_Counter_BTB_N3_10 SAT_Cnt_i_22 ( .SAT_clk(BTB_clk), .SAT_reset(n334), 
        .SAT_enable(n320), .SAT_Ud(n27), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[22]), .SAT_setToDef(s_regenabl_sat[9]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[22]) );
  SAT_Counter_BTB_N3_9 SAT_Cnt_i_23 ( .SAT_clk(BTB_clk), .SAT_reset(n334), 
        .SAT_enable(n319), .SAT_Ud(n27), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[23]), .SAT_setToDef(s_regenabl_sat[8]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[23]) );
  SAT_Counter_BTB_N3_8 SAT_Cnt_i_24 ( .SAT_clk(BTB_clk), .SAT_reset(n334), 
        .SAT_enable(n8), .SAT_Ud(n27), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[24]), .SAT_setToDef(s_regenabl_sat[7]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[24]) );
  SAT_Counter_BTB_N3_7 SAT_Cnt_i_25 ( .SAT_clk(BTB_clk), .SAT_reset(n333), 
        .SAT_enable(n319), .SAT_Ud(n27), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[25]), .SAT_setToDef(s_regenabl_sat[6]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[25]) );
  SAT_Counter_BTB_N3_6 SAT_Cnt_i_26 ( .SAT_clk(BTB_clk), .SAT_reset(n333), 
        .SAT_enable(n320), .SAT_Ud(n27), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[26]), .SAT_setToDef(s_regenabl_sat[5]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[26]) );
  SAT_Counter_BTB_N3_5 SAT_Cnt_i_27 ( .SAT_clk(BTB_clk), .SAT_reset(n333), 
        .SAT_enable(n323), .SAT_Ud(n27), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[27]), .SAT_setToDef(s_regenabl_sat[4]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[27]) );
  SAT_Counter_BTB_N3_4 SAT_Cnt_i_28 ( .SAT_clk(BTB_clk), .SAT_reset(n333), 
        .SAT_enable(n8), .SAT_Ud(n27), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[28]), .SAT_setToDef(s_regenabl_sat[3]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[28]) );
  SAT_Counter_BTB_N3_3 SAT_Cnt_i_29 ( .SAT_clk(BTB_clk), .SAT_reset(n333), 
        .SAT_enable(n318), .SAT_Ud(n27), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[29]), .SAT_setToDef(s_regenabl_sat[2]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[29]) );
  SAT_Counter_BTB_N3_2 SAT_Cnt_i_30 ( .SAT_clk(BTB_clk), .SAT_reset(n333), 
        .SAT_enable(n321), .SAT_Ud(n27), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[30]), .SAT_setToDef(s_regenabl_sat[1]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[30]) );
  SAT_Counter_BTB_N3_1 SAT_Cnt_i_31 ( .SAT_clk(BTB_clk), .SAT_reset(n333), 
        .SAT_enable(n318), .SAT_Ud(n27), .SAT_update(
        s_updateSat_FregCmpBits_Tsats[31]), .SAT_setToDef(s_regenabl_sat[0]), 
        .SAT_SO(s_prediction_Fsat_Tmuxes[31]) );
  Mux_Bit_NBIT_Sel5 MuxSat ( .inputs(s_prediction_Fsat_Tmuxes), .sel({
        s_selmuxes_Fencoder_Tmuxes[4:3], n26, n25, n11}), .\output (
        s_sat_prediction_Toutput) );
  Mux_1Bit_2X1_5 MuxSatOut ( .port0(1'b0), .port1(s_sat_prediction_Toutput), 
        .sel(s_HIT_miss), .portY(s_btb_prediction) );
  Mux_1Bit_2X1_4 Mux_restore ( .port0(s_btb_prediction), .port1(n29), .sel(
        BTB_restore), .portY(BTB_prediction) );
  Mux_NBit_2x1_NBIT_IN32_121 MUX1_0_0 ( .port0({\s_mux_signals[0][0][31] , 
        \s_mux_signals[0][0][30] , \s_mux_signals[0][0][29] , 
        \s_mux_signals[0][0][28] , \s_mux_signals[0][0][27] , 
        \s_mux_signals[0][0][26] , \s_mux_signals[0][0][25] , 
        \s_mux_signals[0][0][24] , \s_mux_signals[0][0][23] , 
        \s_mux_signals[0][0][22] , \s_mux_signals[0][0][21] , 
        \s_mux_signals[0][0][20] , \s_mux_signals[0][0][19] , 
        \s_mux_signals[0][0][18] , \s_mux_signals[0][0][17] , 
        \s_mux_signals[0][0][16] , \s_mux_signals[0][0][15] , 
        \s_mux_signals[0][0][14] , \s_mux_signals[0][0][13] , 
        \s_mux_signals[0][0][12] , \s_mux_signals[0][0][11] , 
        \s_mux_signals[0][0][10] , \s_mux_signals[0][0][9] , 
        \s_mux_signals[0][0][8] , \s_mux_signals[0][0][7] , 
        \s_mux_signals[0][0][6] , \s_mux_signals[0][0][5] , 
        \s_mux_signals[0][0][4] , \s_mux_signals[0][0][3] , 
        \s_mux_signals[0][0][2] , \s_mux_signals[0][0][1] , 
        \s_mux_signals[0][0][0] }), .port1({\s_mux_signals[0][1][31] , 
        \s_mux_signals[0][1][30] , \s_mux_signals[0][1][29] , 
        \s_mux_signals[0][1][28] , \s_mux_signals[0][1][27] , 
        \s_mux_signals[0][1][26] , \s_mux_signals[0][1][25] , 
        \s_mux_signals[0][1][24] , \s_mux_signals[0][1][23] , 
        \s_mux_signals[0][1][22] , \s_mux_signals[0][1][21] , 
        \s_mux_signals[0][1][20] , \s_mux_signals[0][1][19] , 
        \s_mux_signals[0][1][18] , \s_mux_signals[0][1][17] , 
        \s_mux_signals[0][1][16] , \s_mux_signals[0][1][15] , 
        \s_mux_signals[0][1][14] , \s_mux_signals[0][1][13] , 
        \s_mux_signals[0][1][12] , \s_mux_signals[0][1][11] , 
        \s_mux_signals[0][1][10] , \s_mux_signals[0][1][9] , 
        \s_mux_signals[0][1][8] , \s_mux_signals[0][1][7] , 
        \s_mux_signals[0][1][6] , \s_mux_signals[0][1][5] , 
        \s_mux_signals[0][1][4] , \s_mux_signals[0][1][3] , 
        \s_mux_signals[0][1][2] , \s_mux_signals[0][1][1] , 
        \s_mux_signals[0][1][0] }), .sel(n13), .portY({
        \s_mux_signals[1][0][31] , \s_mux_signals[1][0][30] , 
        \s_mux_signals[1][0][29] , \s_mux_signals[1][0][28] , 
        \s_mux_signals[1][0][27] , \s_mux_signals[1][0][26] , 
        \s_mux_signals[1][0][25] , \s_mux_signals[1][0][24] , 
        \s_mux_signals[1][0][23] , \s_mux_signals[1][0][22] , 
        \s_mux_signals[1][0][21] , \s_mux_signals[1][0][20] , 
        \s_mux_signals[1][0][19] , \s_mux_signals[1][0][18] , 
        \s_mux_signals[1][0][17] , \s_mux_signals[1][0][16] , 
        \s_mux_signals[1][0][15] , \s_mux_signals[1][0][14] , 
        \s_mux_signals[1][0][13] , \s_mux_signals[1][0][12] , 
        \s_mux_signals[1][0][11] , \s_mux_signals[1][0][10] , 
        \s_mux_signals[1][0][9] , \s_mux_signals[1][0][8] , 
        \s_mux_signals[1][0][7] , \s_mux_signals[1][0][6] , 
        \s_mux_signals[1][0][5] , \s_mux_signals[1][0][4] , 
        \s_mux_signals[1][0][3] , \s_mux_signals[1][0][2] , 
        \s_mux_signals[1][0][1] , \s_mux_signals[1][0][0] }) );
  Mux_NBit_2x1_NBIT_IN32_120 MUX1_0_2 ( .port0({\s_mux_signals[0][2][31] , 
        \s_mux_signals[0][2][30] , \s_mux_signals[0][2][29] , 
        \s_mux_signals[0][2][28] , \s_mux_signals[0][2][27] , 
        \s_mux_signals[0][2][26] , \s_mux_signals[0][2][25] , 
        \s_mux_signals[0][2][24] , \s_mux_signals[0][2][23] , 
        \s_mux_signals[0][2][22] , \s_mux_signals[0][2][21] , 
        \s_mux_signals[0][2][20] , \s_mux_signals[0][2][19] , 
        \s_mux_signals[0][2][18] , \s_mux_signals[0][2][17] , 
        \s_mux_signals[0][2][16] , \s_mux_signals[0][2][15] , 
        \s_mux_signals[0][2][14] , \s_mux_signals[0][2][13] , 
        \s_mux_signals[0][2][12] , \s_mux_signals[0][2][11] , 
        \s_mux_signals[0][2][10] , \s_mux_signals[0][2][9] , 
        \s_mux_signals[0][2][8] , \s_mux_signals[0][2][7] , 
        \s_mux_signals[0][2][6] , \s_mux_signals[0][2][5] , 
        \s_mux_signals[0][2][4] , \s_mux_signals[0][2][3] , 
        \s_mux_signals[0][2][2] , \s_mux_signals[0][2][1] , 
        \s_mux_signals[0][2][0] }), .port1({\s_mux_signals[0][3][31] , 
        \s_mux_signals[0][3][30] , \s_mux_signals[0][3][29] , 
        \s_mux_signals[0][3][28] , \s_mux_signals[0][3][27] , 
        \s_mux_signals[0][3][26] , \s_mux_signals[0][3][25] , 
        \s_mux_signals[0][3][24] , \s_mux_signals[0][3][23] , 
        \s_mux_signals[0][3][22] , \s_mux_signals[0][3][21] , 
        \s_mux_signals[0][3][20] , \s_mux_signals[0][3][19] , 
        \s_mux_signals[0][3][18] , \s_mux_signals[0][3][17] , 
        \s_mux_signals[0][3][16] , \s_mux_signals[0][3][15] , 
        \s_mux_signals[0][3][14] , \s_mux_signals[0][3][13] , 
        \s_mux_signals[0][3][12] , \s_mux_signals[0][3][11] , 
        \s_mux_signals[0][3][10] , \s_mux_signals[0][3][9] , 
        \s_mux_signals[0][3][8] , \s_mux_signals[0][3][7] , 
        \s_mux_signals[0][3][6] , \s_mux_signals[0][3][5] , 
        \s_mux_signals[0][3][4] , \s_mux_signals[0][3][3] , 
        \s_mux_signals[0][3][2] , \s_mux_signals[0][3][1] , 
        \s_mux_signals[0][3][0] }), .sel(n11), .portY({
        \s_mux_signals[1][2][31] , \s_mux_signals[1][2][30] , 
        \s_mux_signals[1][2][29] , \s_mux_signals[1][2][28] , 
        \s_mux_signals[1][2][27] , \s_mux_signals[1][2][26] , 
        \s_mux_signals[1][2][25] , \s_mux_signals[1][2][24] , 
        \s_mux_signals[1][2][23] , \s_mux_signals[1][2][22] , 
        \s_mux_signals[1][2][21] , \s_mux_signals[1][2][20] , 
        \s_mux_signals[1][2][19] , \s_mux_signals[1][2][18] , 
        \s_mux_signals[1][2][17] , \s_mux_signals[1][2][16] , 
        \s_mux_signals[1][2][15] , \s_mux_signals[1][2][14] , 
        \s_mux_signals[1][2][13] , \s_mux_signals[1][2][12] , 
        \s_mux_signals[1][2][11] , \s_mux_signals[1][2][10] , 
        \s_mux_signals[1][2][9] , \s_mux_signals[1][2][8] , 
        \s_mux_signals[1][2][7] , \s_mux_signals[1][2][6] , 
        \s_mux_signals[1][2][5] , \s_mux_signals[1][2][4] , 
        \s_mux_signals[1][2][3] , \s_mux_signals[1][2][2] , 
        \s_mux_signals[1][2][1] , \s_mux_signals[1][2][0] }) );
  Mux_NBit_2x1_NBIT_IN32_119 MUX1_0_4 ( .port0({\s_mux_signals[0][4][31] , 
        \s_mux_signals[0][4][30] , \s_mux_signals[0][4][29] , 
        \s_mux_signals[0][4][28] , \s_mux_signals[0][4][27] , 
        \s_mux_signals[0][4][26] , \s_mux_signals[0][4][25] , 
        \s_mux_signals[0][4][24] , \s_mux_signals[0][4][23] , 
        \s_mux_signals[0][4][22] , \s_mux_signals[0][4][21] , 
        \s_mux_signals[0][4][20] , \s_mux_signals[0][4][19] , 
        \s_mux_signals[0][4][18] , \s_mux_signals[0][4][17] , 
        \s_mux_signals[0][4][16] , \s_mux_signals[0][4][15] , 
        \s_mux_signals[0][4][14] , \s_mux_signals[0][4][13] , 
        \s_mux_signals[0][4][12] , \s_mux_signals[0][4][11] , 
        \s_mux_signals[0][4][10] , \s_mux_signals[0][4][9] , 
        \s_mux_signals[0][4][8] , \s_mux_signals[0][4][7] , 
        \s_mux_signals[0][4][6] , \s_mux_signals[0][4][5] , 
        \s_mux_signals[0][4][4] , \s_mux_signals[0][4][3] , 
        \s_mux_signals[0][4][2] , \s_mux_signals[0][4][1] , 
        \s_mux_signals[0][4][0] }), .port1({\s_mux_signals[0][5][31] , 
        \s_mux_signals[0][5][30] , \s_mux_signals[0][5][29] , 
        \s_mux_signals[0][5][28] , \s_mux_signals[0][5][27] , 
        \s_mux_signals[0][5][26] , \s_mux_signals[0][5][25] , 
        \s_mux_signals[0][5][24] , \s_mux_signals[0][5][23] , 
        \s_mux_signals[0][5][22] , \s_mux_signals[0][5][21] , 
        \s_mux_signals[0][5][20] , \s_mux_signals[0][5][19] , 
        \s_mux_signals[0][5][18] , \s_mux_signals[0][5][17] , 
        \s_mux_signals[0][5][16] , \s_mux_signals[0][5][15] , 
        \s_mux_signals[0][5][14] , \s_mux_signals[0][5][13] , 
        \s_mux_signals[0][5][12] , \s_mux_signals[0][5][11] , 
        \s_mux_signals[0][5][10] , \s_mux_signals[0][5][9] , 
        \s_mux_signals[0][5][8] , \s_mux_signals[0][5][7] , 
        \s_mux_signals[0][5][6] , \s_mux_signals[0][5][5] , 
        \s_mux_signals[0][5][4] , \s_mux_signals[0][5][3] , 
        \s_mux_signals[0][5][2] , \s_mux_signals[0][5][1] , 
        \s_mux_signals[0][5][0] }), .sel(n11), .portY({
        \s_mux_signals[1][4][31] , \s_mux_signals[1][4][30] , 
        \s_mux_signals[1][4][29] , \s_mux_signals[1][4][28] , 
        \s_mux_signals[1][4][27] , \s_mux_signals[1][4][26] , 
        \s_mux_signals[1][4][25] , \s_mux_signals[1][4][24] , 
        \s_mux_signals[1][4][23] , \s_mux_signals[1][4][22] , 
        \s_mux_signals[1][4][21] , \s_mux_signals[1][4][20] , 
        \s_mux_signals[1][4][19] , \s_mux_signals[1][4][18] , 
        \s_mux_signals[1][4][17] , \s_mux_signals[1][4][16] , 
        \s_mux_signals[1][4][15] , \s_mux_signals[1][4][14] , 
        \s_mux_signals[1][4][13] , \s_mux_signals[1][4][12] , 
        \s_mux_signals[1][4][11] , \s_mux_signals[1][4][10] , 
        \s_mux_signals[1][4][9] , \s_mux_signals[1][4][8] , 
        \s_mux_signals[1][4][7] , \s_mux_signals[1][4][6] , 
        \s_mux_signals[1][4][5] , \s_mux_signals[1][4][4] , 
        \s_mux_signals[1][4][3] , \s_mux_signals[1][4][2] , 
        \s_mux_signals[1][4][1] , \s_mux_signals[1][4][0] }) );
  Mux_NBit_2x1_NBIT_IN32_118 MUX1_0_6 ( .port0({\s_mux_signals[0][6][31] , 
        \s_mux_signals[0][6][30] , \s_mux_signals[0][6][29] , 
        \s_mux_signals[0][6][28] , \s_mux_signals[0][6][27] , 
        \s_mux_signals[0][6][26] , \s_mux_signals[0][6][25] , 
        \s_mux_signals[0][6][24] , \s_mux_signals[0][6][23] , 
        \s_mux_signals[0][6][22] , \s_mux_signals[0][6][21] , 
        \s_mux_signals[0][6][20] , \s_mux_signals[0][6][19] , 
        \s_mux_signals[0][6][18] , \s_mux_signals[0][6][17] , 
        \s_mux_signals[0][6][16] , \s_mux_signals[0][6][15] , 
        \s_mux_signals[0][6][14] , \s_mux_signals[0][6][13] , 
        \s_mux_signals[0][6][12] , \s_mux_signals[0][6][11] , 
        \s_mux_signals[0][6][10] , \s_mux_signals[0][6][9] , 
        \s_mux_signals[0][6][8] , \s_mux_signals[0][6][7] , 
        \s_mux_signals[0][6][6] , \s_mux_signals[0][6][5] , 
        \s_mux_signals[0][6][4] , \s_mux_signals[0][6][3] , 
        \s_mux_signals[0][6][2] , \s_mux_signals[0][6][1] , 
        \s_mux_signals[0][6][0] }), .port1({\s_mux_signals[0][7][31] , 
        \s_mux_signals[0][7][30] , \s_mux_signals[0][7][29] , 
        \s_mux_signals[0][7][28] , \s_mux_signals[0][7][27] , 
        \s_mux_signals[0][7][26] , \s_mux_signals[0][7][25] , 
        \s_mux_signals[0][7][24] , \s_mux_signals[0][7][23] , 
        \s_mux_signals[0][7][22] , \s_mux_signals[0][7][21] , 
        \s_mux_signals[0][7][20] , \s_mux_signals[0][7][19] , 
        \s_mux_signals[0][7][18] , \s_mux_signals[0][7][17] , 
        \s_mux_signals[0][7][16] , \s_mux_signals[0][7][15] , 
        \s_mux_signals[0][7][14] , \s_mux_signals[0][7][13] , 
        \s_mux_signals[0][7][12] , \s_mux_signals[0][7][11] , 
        \s_mux_signals[0][7][10] , \s_mux_signals[0][7][9] , 
        \s_mux_signals[0][7][8] , \s_mux_signals[0][7][7] , 
        \s_mux_signals[0][7][6] , \s_mux_signals[0][7][5] , 
        \s_mux_signals[0][7][4] , \s_mux_signals[0][7][3] , 
        \s_mux_signals[0][7][2] , \s_mux_signals[0][7][1] , 
        \s_mux_signals[0][7][0] }), .sel(n11), .portY({
        \s_mux_signals[1][6][31] , \s_mux_signals[1][6][30] , 
        \s_mux_signals[1][6][29] , \s_mux_signals[1][6][28] , 
        \s_mux_signals[1][6][27] , \s_mux_signals[1][6][26] , 
        \s_mux_signals[1][6][25] , \s_mux_signals[1][6][24] , 
        \s_mux_signals[1][6][23] , \s_mux_signals[1][6][22] , 
        \s_mux_signals[1][6][21] , \s_mux_signals[1][6][20] , 
        \s_mux_signals[1][6][19] , \s_mux_signals[1][6][18] , 
        \s_mux_signals[1][6][17] , \s_mux_signals[1][6][16] , 
        \s_mux_signals[1][6][15] , \s_mux_signals[1][6][14] , 
        \s_mux_signals[1][6][13] , \s_mux_signals[1][6][12] , 
        \s_mux_signals[1][6][11] , \s_mux_signals[1][6][10] , 
        \s_mux_signals[1][6][9] , \s_mux_signals[1][6][8] , 
        \s_mux_signals[1][6][7] , \s_mux_signals[1][6][6] , 
        \s_mux_signals[1][6][5] , \s_mux_signals[1][6][4] , 
        \s_mux_signals[1][6][3] , \s_mux_signals[1][6][2] , 
        \s_mux_signals[1][6][1] , \s_mux_signals[1][6][0] }) );
  Mux_NBit_2x1_NBIT_IN32_117 MUX1_0_8 ( .port0({\s_mux_signals[0][8][31] , 
        \s_mux_signals[0][8][30] , \s_mux_signals[0][8][29] , 
        \s_mux_signals[0][8][28] , \s_mux_signals[0][8][27] , 
        \s_mux_signals[0][8][26] , \s_mux_signals[0][8][25] , 
        \s_mux_signals[0][8][24] , \s_mux_signals[0][8][23] , 
        \s_mux_signals[0][8][22] , \s_mux_signals[0][8][21] , 
        \s_mux_signals[0][8][20] , \s_mux_signals[0][8][19] , 
        \s_mux_signals[0][8][18] , \s_mux_signals[0][8][17] , 
        \s_mux_signals[0][8][16] , \s_mux_signals[0][8][15] , 
        \s_mux_signals[0][8][14] , \s_mux_signals[0][8][13] , 
        \s_mux_signals[0][8][12] , \s_mux_signals[0][8][11] , 
        \s_mux_signals[0][8][10] , \s_mux_signals[0][8][9] , 
        \s_mux_signals[0][8][8] , \s_mux_signals[0][8][7] , 
        \s_mux_signals[0][8][6] , \s_mux_signals[0][8][5] , 
        \s_mux_signals[0][8][4] , \s_mux_signals[0][8][3] , 
        \s_mux_signals[0][8][2] , \s_mux_signals[0][8][1] , 
        \s_mux_signals[0][8][0] }), .port1({\s_mux_signals[0][9][31] , 
        \s_mux_signals[0][9][30] , \s_mux_signals[0][9][29] , 
        \s_mux_signals[0][9][28] , \s_mux_signals[0][9][27] , 
        \s_mux_signals[0][9][26] , \s_mux_signals[0][9][25] , 
        \s_mux_signals[0][9][24] , \s_mux_signals[0][9][23] , 
        \s_mux_signals[0][9][22] , \s_mux_signals[0][9][21] , 
        \s_mux_signals[0][9][20] , \s_mux_signals[0][9][19] , 
        \s_mux_signals[0][9][18] , \s_mux_signals[0][9][17] , 
        \s_mux_signals[0][9][16] , \s_mux_signals[0][9][15] , 
        \s_mux_signals[0][9][14] , \s_mux_signals[0][9][13] , 
        \s_mux_signals[0][9][12] , \s_mux_signals[0][9][11] , 
        \s_mux_signals[0][9][10] , \s_mux_signals[0][9][9] , 
        \s_mux_signals[0][9][8] , \s_mux_signals[0][9][7] , 
        \s_mux_signals[0][9][6] , \s_mux_signals[0][9][5] , 
        \s_mux_signals[0][9][4] , \s_mux_signals[0][9][3] , 
        \s_mux_signals[0][9][2] , \s_mux_signals[0][9][1] , 
        \s_mux_signals[0][9][0] }), .sel(n11), .portY({
        \s_mux_signals[1][8][31] , \s_mux_signals[1][8][30] , 
        \s_mux_signals[1][8][29] , \s_mux_signals[1][8][28] , 
        \s_mux_signals[1][8][27] , \s_mux_signals[1][8][26] , 
        \s_mux_signals[1][8][25] , \s_mux_signals[1][8][24] , 
        \s_mux_signals[1][8][23] , \s_mux_signals[1][8][22] , 
        \s_mux_signals[1][8][21] , \s_mux_signals[1][8][20] , 
        \s_mux_signals[1][8][19] , \s_mux_signals[1][8][18] , 
        \s_mux_signals[1][8][17] , \s_mux_signals[1][8][16] , 
        \s_mux_signals[1][8][15] , \s_mux_signals[1][8][14] , 
        \s_mux_signals[1][8][13] , \s_mux_signals[1][8][12] , 
        \s_mux_signals[1][8][11] , \s_mux_signals[1][8][10] , 
        \s_mux_signals[1][8][9] , \s_mux_signals[1][8][8] , 
        \s_mux_signals[1][8][7] , \s_mux_signals[1][8][6] , 
        \s_mux_signals[1][8][5] , \s_mux_signals[1][8][4] , 
        \s_mux_signals[1][8][3] , \s_mux_signals[1][8][2] , 
        \s_mux_signals[1][8][1] , \s_mux_signals[1][8][0] }) );
  Mux_NBit_2x1_NBIT_IN32_116 MUX1_0_10 ( .port0({\s_mux_signals[0][10][31] , 
        \s_mux_signals[0][10][30] , \s_mux_signals[0][10][29] , 
        \s_mux_signals[0][10][28] , \s_mux_signals[0][10][27] , 
        \s_mux_signals[0][10][26] , \s_mux_signals[0][10][25] , 
        \s_mux_signals[0][10][24] , \s_mux_signals[0][10][23] , 
        \s_mux_signals[0][10][22] , \s_mux_signals[0][10][21] , 
        \s_mux_signals[0][10][20] , \s_mux_signals[0][10][19] , 
        \s_mux_signals[0][10][18] , \s_mux_signals[0][10][17] , 
        \s_mux_signals[0][10][16] , \s_mux_signals[0][10][15] , 
        \s_mux_signals[0][10][14] , \s_mux_signals[0][10][13] , 
        \s_mux_signals[0][10][12] , \s_mux_signals[0][10][11] , 
        \s_mux_signals[0][10][10] , \s_mux_signals[0][10][9] , 
        \s_mux_signals[0][10][8] , \s_mux_signals[0][10][7] , 
        \s_mux_signals[0][10][6] , \s_mux_signals[0][10][5] , 
        \s_mux_signals[0][10][4] , \s_mux_signals[0][10][3] , 
        \s_mux_signals[0][10][2] , \s_mux_signals[0][10][1] , 
        \s_mux_signals[0][10][0] }), .port1({\s_mux_signals[0][11][31] , 
        \s_mux_signals[0][11][30] , \s_mux_signals[0][11][29] , 
        \s_mux_signals[0][11][28] , \s_mux_signals[0][11][27] , 
        \s_mux_signals[0][11][26] , \s_mux_signals[0][11][25] , 
        \s_mux_signals[0][11][24] , \s_mux_signals[0][11][23] , 
        \s_mux_signals[0][11][22] , \s_mux_signals[0][11][21] , 
        \s_mux_signals[0][11][20] , \s_mux_signals[0][11][19] , 
        \s_mux_signals[0][11][18] , \s_mux_signals[0][11][17] , 
        \s_mux_signals[0][11][16] , \s_mux_signals[0][11][15] , 
        \s_mux_signals[0][11][14] , \s_mux_signals[0][11][13] , 
        \s_mux_signals[0][11][12] , \s_mux_signals[0][11][11] , 
        \s_mux_signals[0][11][10] , \s_mux_signals[0][11][9] , 
        \s_mux_signals[0][11][8] , \s_mux_signals[0][11][7] , 
        \s_mux_signals[0][11][6] , \s_mux_signals[0][11][5] , 
        \s_mux_signals[0][11][4] , \s_mux_signals[0][11][3] , 
        \s_mux_signals[0][11][2] , \s_mux_signals[0][11][1] , 
        \s_mux_signals[0][11][0] }), .sel(n11), .portY({
        \s_mux_signals[1][10][31] , \s_mux_signals[1][10][30] , 
        \s_mux_signals[1][10][29] , \s_mux_signals[1][10][28] , 
        \s_mux_signals[1][10][27] , \s_mux_signals[1][10][26] , 
        \s_mux_signals[1][10][25] , \s_mux_signals[1][10][24] , 
        \s_mux_signals[1][10][23] , \s_mux_signals[1][10][22] , 
        \s_mux_signals[1][10][21] , \s_mux_signals[1][10][20] , 
        \s_mux_signals[1][10][19] , \s_mux_signals[1][10][18] , 
        \s_mux_signals[1][10][17] , \s_mux_signals[1][10][16] , 
        \s_mux_signals[1][10][15] , \s_mux_signals[1][10][14] , 
        \s_mux_signals[1][10][13] , \s_mux_signals[1][10][12] , 
        \s_mux_signals[1][10][11] , \s_mux_signals[1][10][10] , 
        \s_mux_signals[1][10][9] , \s_mux_signals[1][10][8] , 
        \s_mux_signals[1][10][7] , \s_mux_signals[1][10][6] , 
        \s_mux_signals[1][10][5] , \s_mux_signals[1][10][4] , 
        \s_mux_signals[1][10][3] , \s_mux_signals[1][10][2] , 
        \s_mux_signals[1][10][1] , \s_mux_signals[1][10][0] }) );
  Mux_NBit_2x1_NBIT_IN32_115 MUX1_0_12 ( .port0({\s_mux_signals[0][12][31] , 
        \s_mux_signals[0][12][30] , \s_mux_signals[0][12][29] , 
        \s_mux_signals[0][12][28] , \s_mux_signals[0][12][27] , 
        \s_mux_signals[0][12][26] , \s_mux_signals[0][12][25] , 
        \s_mux_signals[0][12][24] , \s_mux_signals[0][12][23] , 
        \s_mux_signals[0][12][22] , \s_mux_signals[0][12][21] , 
        \s_mux_signals[0][12][20] , \s_mux_signals[0][12][19] , 
        \s_mux_signals[0][12][18] , \s_mux_signals[0][12][17] , 
        \s_mux_signals[0][12][16] , \s_mux_signals[0][12][15] , 
        \s_mux_signals[0][12][14] , \s_mux_signals[0][12][13] , 
        \s_mux_signals[0][12][12] , \s_mux_signals[0][12][11] , 
        \s_mux_signals[0][12][10] , \s_mux_signals[0][12][9] , 
        \s_mux_signals[0][12][8] , \s_mux_signals[0][12][7] , 
        \s_mux_signals[0][12][6] , \s_mux_signals[0][12][5] , 
        \s_mux_signals[0][12][4] , \s_mux_signals[0][12][3] , 
        \s_mux_signals[0][12][2] , \s_mux_signals[0][12][1] , 
        \s_mux_signals[0][12][0] }), .port1({\s_mux_signals[0][13][31] , 
        \s_mux_signals[0][13][30] , \s_mux_signals[0][13][29] , 
        \s_mux_signals[0][13][28] , \s_mux_signals[0][13][27] , 
        \s_mux_signals[0][13][26] , \s_mux_signals[0][13][25] , 
        \s_mux_signals[0][13][24] , \s_mux_signals[0][13][23] , 
        \s_mux_signals[0][13][22] , \s_mux_signals[0][13][21] , 
        \s_mux_signals[0][13][20] , \s_mux_signals[0][13][19] , 
        \s_mux_signals[0][13][18] , \s_mux_signals[0][13][17] , 
        \s_mux_signals[0][13][16] , \s_mux_signals[0][13][15] , 
        \s_mux_signals[0][13][14] , \s_mux_signals[0][13][13] , 
        \s_mux_signals[0][13][12] , \s_mux_signals[0][13][11] , 
        \s_mux_signals[0][13][10] , \s_mux_signals[0][13][9] , 
        \s_mux_signals[0][13][8] , \s_mux_signals[0][13][7] , 
        \s_mux_signals[0][13][6] , \s_mux_signals[0][13][5] , 
        \s_mux_signals[0][13][4] , \s_mux_signals[0][13][3] , 
        \s_mux_signals[0][13][2] , \s_mux_signals[0][13][1] , 
        \s_mux_signals[0][13][0] }), .sel(n11), .portY({
        \s_mux_signals[1][12][31] , \s_mux_signals[1][12][30] , 
        \s_mux_signals[1][12][29] , \s_mux_signals[1][12][28] , 
        \s_mux_signals[1][12][27] , \s_mux_signals[1][12][26] , 
        \s_mux_signals[1][12][25] , \s_mux_signals[1][12][24] , 
        \s_mux_signals[1][12][23] , \s_mux_signals[1][12][22] , 
        \s_mux_signals[1][12][21] , \s_mux_signals[1][12][20] , 
        \s_mux_signals[1][12][19] , \s_mux_signals[1][12][18] , 
        \s_mux_signals[1][12][17] , \s_mux_signals[1][12][16] , 
        \s_mux_signals[1][12][15] , \s_mux_signals[1][12][14] , 
        \s_mux_signals[1][12][13] , \s_mux_signals[1][12][12] , 
        \s_mux_signals[1][12][11] , \s_mux_signals[1][12][10] , 
        \s_mux_signals[1][12][9] , \s_mux_signals[1][12][8] , 
        \s_mux_signals[1][12][7] , \s_mux_signals[1][12][6] , 
        \s_mux_signals[1][12][5] , \s_mux_signals[1][12][4] , 
        \s_mux_signals[1][12][3] , \s_mux_signals[1][12][2] , 
        \s_mux_signals[1][12][1] , \s_mux_signals[1][12][0] }) );
  Mux_NBit_2x1_NBIT_IN32_114 MUX1_0_14 ( .port0({\s_mux_signals[0][14][31] , 
        \s_mux_signals[0][14][30] , \s_mux_signals[0][14][29] , 
        \s_mux_signals[0][14][28] , \s_mux_signals[0][14][27] , 
        \s_mux_signals[0][14][26] , \s_mux_signals[0][14][25] , 
        \s_mux_signals[0][14][24] , \s_mux_signals[0][14][23] , 
        \s_mux_signals[0][14][22] , \s_mux_signals[0][14][21] , 
        \s_mux_signals[0][14][20] , \s_mux_signals[0][14][19] , 
        \s_mux_signals[0][14][18] , \s_mux_signals[0][14][17] , 
        \s_mux_signals[0][14][16] , \s_mux_signals[0][14][15] , 
        \s_mux_signals[0][14][14] , \s_mux_signals[0][14][13] , 
        \s_mux_signals[0][14][12] , \s_mux_signals[0][14][11] , 
        \s_mux_signals[0][14][10] , \s_mux_signals[0][14][9] , 
        \s_mux_signals[0][14][8] , \s_mux_signals[0][14][7] , 
        \s_mux_signals[0][14][6] , \s_mux_signals[0][14][5] , 
        \s_mux_signals[0][14][4] , \s_mux_signals[0][14][3] , 
        \s_mux_signals[0][14][2] , \s_mux_signals[0][14][1] , 
        \s_mux_signals[0][14][0] }), .port1({\s_mux_signals[0][15][31] , 
        \s_mux_signals[0][15][30] , \s_mux_signals[0][15][29] , 
        \s_mux_signals[0][15][28] , \s_mux_signals[0][15][27] , 
        \s_mux_signals[0][15][26] , \s_mux_signals[0][15][25] , 
        \s_mux_signals[0][15][24] , \s_mux_signals[0][15][23] , 
        \s_mux_signals[0][15][22] , \s_mux_signals[0][15][21] , 
        \s_mux_signals[0][15][20] , \s_mux_signals[0][15][19] , 
        \s_mux_signals[0][15][18] , \s_mux_signals[0][15][17] , 
        \s_mux_signals[0][15][16] , \s_mux_signals[0][15][15] , 
        \s_mux_signals[0][15][14] , \s_mux_signals[0][15][13] , 
        \s_mux_signals[0][15][12] , \s_mux_signals[0][15][11] , 
        \s_mux_signals[0][15][10] , \s_mux_signals[0][15][9] , 
        \s_mux_signals[0][15][8] , \s_mux_signals[0][15][7] , 
        \s_mux_signals[0][15][6] , \s_mux_signals[0][15][5] , 
        \s_mux_signals[0][15][4] , \s_mux_signals[0][15][3] , 
        \s_mux_signals[0][15][2] , \s_mux_signals[0][15][1] , 
        \s_mux_signals[0][15][0] }), .sel(n11), .portY({
        \s_mux_signals[1][14][31] , \s_mux_signals[1][14][30] , 
        \s_mux_signals[1][14][29] , \s_mux_signals[1][14][28] , 
        \s_mux_signals[1][14][27] , \s_mux_signals[1][14][26] , 
        \s_mux_signals[1][14][25] , \s_mux_signals[1][14][24] , 
        \s_mux_signals[1][14][23] , \s_mux_signals[1][14][22] , 
        \s_mux_signals[1][14][21] , \s_mux_signals[1][14][20] , 
        \s_mux_signals[1][14][19] , \s_mux_signals[1][14][18] , 
        \s_mux_signals[1][14][17] , \s_mux_signals[1][14][16] , 
        \s_mux_signals[1][14][15] , \s_mux_signals[1][14][14] , 
        \s_mux_signals[1][14][13] , \s_mux_signals[1][14][12] , 
        \s_mux_signals[1][14][11] , \s_mux_signals[1][14][10] , 
        \s_mux_signals[1][14][9] , \s_mux_signals[1][14][8] , 
        \s_mux_signals[1][14][7] , \s_mux_signals[1][14][6] , 
        \s_mux_signals[1][14][5] , \s_mux_signals[1][14][4] , 
        \s_mux_signals[1][14][3] , \s_mux_signals[1][14][2] , 
        \s_mux_signals[1][14][1] , \s_mux_signals[1][14][0] }) );
  Mux_NBit_2x1_NBIT_IN32_113 MUX1_0_16 ( .port0({\s_mux_signals[0][16][31] , 
        \s_mux_signals[0][16][30] , \s_mux_signals[0][16][29] , 
        \s_mux_signals[0][16][28] , \s_mux_signals[0][16][27] , 
        \s_mux_signals[0][16][26] , \s_mux_signals[0][16][25] , 
        \s_mux_signals[0][16][24] , \s_mux_signals[0][16][23] , 
        \s_mux_signals[0][16][22] , \s_mux_signals[0][16][21] , 
        \s_mux_signals[0][16][20] , \s_mux_signals[0][16][19] , 
        \s_mux_signals[0][16][18] , \s_mux_signals[0][16][17] , 
        \s_mux_signals[0][16][16] , \s_mux_signals[0][16][15] , 
        \s_mux_signals[0][16][14] , \s_mux_signals[0][16][13] , 
        \s_mux_signals[0][16][12] , \s_mux_signals[0][16][11] , 
        \s_mux_signals[0][16][10] , \s_mux_signals[0][16][9] , 
        \s_mux_signals[0][16][8] , \s_mux_signals[0][16][7] , 
        \s_mux_signals[0][16][6] , \s_mux_signals[0][16][5] , 
        \s_mux_signals[0][16][4] , \s_mux_signals[0][16][3] , 
        \s_mux_signals[0][16][2] , \s_mux_signals[0][16][1] , 
        \s_mux_signals[0][16][0] }), .port1({\s_mux_signals[0][17][31] , 
        \s_mux_signals[0][17][30] , \s_mux_signals[0][17][29] , 
        \s_mux_signals[0][17][28] , \s_mux_signals[0][17][27] , 
        \s_mux_signals[0][17][26] , \s_mux_signals[0][17][25] , 
        \s_mux_signals[0][17][24] , \s_mux_signals[0][17][23] , 
        \s_mux_signals[0][17][22] , \s_mux_signals[0][17][21] , 
        \s_mux_signals[0][17][20] , \s_mux_signals[0][17][19] , 
        \s_mux_signals[0][17][18] , \s_mux_signals[0][17][17] , 
        \s_mux_signals[0][17][16] , \s_mux_signals[0][17][15] , 
        \s_mux_signals[0][17][14] , \s_mux_signals[0][17][13] , 
        \s_mux_signals[0][17][12] , \s_mux_signals[0][17][11] , 
        \s_mux_signals[0][17][10] , \s_mux_signals[0][17][9] , 
        \s_mux_signals[0][17][8] , \s_mux_signals[0][17][7] , 
        \s_mux_signals[0][17][6] , \s_mux_signals[0][17][5] , 
        \s_mux_signals[0][17][4] , \s_mux_signals[0][17][3] , 
        \s_mux_signals[0][17][2] , \s_mux_signals[0][17][1] , 
        \s_mux_signals[0][17][0] }), .sel(n12), .portY({
        \s_mux_signals[1][16][31] , \s_mux_signals[1][16][30] , 
        \s_mux_signals[1][16][29] , \s_mux_signals[1][16][28] , 
        \s_mux_signals[1][16][27] , \s_mux_signals[1][16][26] , 
        \s_mux_signals[1][16][25] , \s_mux_signals[1][16][24] , 
        \s_mux_signals[1][16][23] , \s_mux_signals[1][16][22] , 
        \s_mux_signals[1][16][21] , \s_mux_signals[1][16][20] , 
        \s_mux_signals[1][16][19] , \s_mux_signals[1][16][18] , 
        \s_mux_signals[1][16][17] , \s_mux_signals[1][16][16] , 
        \s_mux_signals[1][16][15] , \s_mux_signals[1][16][14] , 
        \s_mux_signals[1][16][13] , \s_mux_signals[1][16][12] , 
        \s_mux_signals[1][16][11] , \s_mux_signals[1][16][10] , 
        \s_mux_signals[1][16][9] , \s_mux_signals[1][16][8] , 
        \s_mux_signals[1][16][7] , \s_mux_signals[1][16][6] , 
        \s_mux_signals[1][16][5] , \s_mux_signals[1][16][4] , 
        \s_mux_signals[1][16][3] , \s_mux_signals[1][16][2] , 
        \s_mux_signals[1][16][1] , \s_mux_signals[1][16][0] }) );
  Mux_NBit_2x1_NBIT_IN32_112 MUX1_0_18 ( .port0({\s_mux_signals[0][18][31] , 
        \s_mux_signals[0][18][30] , \s_mux_signals[0][18][29] , 
        \s_mux_signals[0][18][28] , \s_mux_signals[0][18][27] , 
        \s_mux_signals[0][18][26] , \s_mux_signals[0][18][25] , 
        \s_mux_signals[0][18][24] , \s_mux_signals[0][18][23] , 
        \s_mux_signals[0][18][22] , \s_mux_signals[0][18][21] , 
        \s_mux_signals[0][18][20] , \s_mux_signals[0][18][19] , 
        \s_mux_signals[0][18][18] , \s_mux_signals[0][18][17] , 
        \s_mux_signals[0][18][16] , \s_mux_signals[0][18][15] , 
        \s_mux_signals[0][18][14] , \s_mux_signals[0][18][13] , 
        \s_mux_signals[0][18][12] , \s_mux_signals[0][18][11] , 
        \s_mux_signals[0][18][10] , \s_mux_signals[0][18][9] , 
        \s_mux_signals[0][18][8] , \s_mux_signals[0][18][7] , 
        \s_mux_signals[0][18][6] , \s_mux_signals[0][18][5] , 
        \s_mux_signals[0][18][4] , \s_mux_signals[0][18][3] , 
        \s_mux_signals[0][18][2] , \s_mux_signals[0][18][1] , 
        \s_mux_signals[0][18][0] }), .port1({\s_mux_signals[0][19][31] , 
        \s_mux_signals[0][19][30] , \s_mux_signals[0][19][29] , 
        \s_mux_signals[0][19][28] , \s_mux_signals[0][19][27] , 
        \s_mux_signals[0][19][26] , \s_mux_signals[0][19][25] , 
        \s_mux_signals[0][19][24] , \s_mux_signals[0][19][23] , 
        \s_mux_signals[0][19][22] , \s_mux_signals[0][19][21] , 
        \s_mux_signals[0][19][20] , \s_mux_signals[0][19][19] , 
        \s_mux_signals[0][19][18] , \s_mux_signals[0][19][17] , 
        \s_mux_signals[0][19][16] , \s_mux_signals[0][19][15] , 
        \s_mux_signals[0][19][14] , \s_mux_signals[0][19][13] , 
        \s_mux_signals[0][19][12] , \s_mux_signals[0][19][11] , 
        \s_mux_signals[0][19][10] , \s_mux_signals[0][19][9] , 
        \s_mux_signals[0][19][8] , \s_mux_signals[0][19][7] , 
        \s_mux_signals[0][19][6] , \s_mux_signals[0][19][5] , 
        \s_mux_signals[0][19][4] , \s_mux_signals[0][19][3] , 
        \s_mux_signals[0][19][2] , \s_mux_signals[0][19][1] , 
        \s_mux_signals[0][19][0] }), .sel(n12), .portY({
        \s_mux_signals[1][18][31] , \s_mux_signals[1][18][30] , 
        \s_mux_signals[1][18][29] , \s_mux_signals[1][18][28] , 
        \s_mux_signals[1][18][27] , \s_mux_signals[1][18][26] , 
        \s_mux_signals[1][18][25] , \s_mux_signals[1][18][24] , 
        \s_mux_signals[1][18][23] , \s_mux_signals[1][18][22] , 
        \s_mux_signals[1][18][21] , \s_mux_signals[1][18][20] , 
        \s_mux_signals[1][18][19] , \s_mux_signals[1][18][18] , 
        \s_mux_signals[1][18][17] , \s_mux_signals[1][18][16] , 
        \s_mux_signals[1][18][15] , \s_mux_signals[1][18][14] , 
        \s_mux_signals[1][18][13] , \s_mux_signals[1][18][12] , 
        \s_mux_signals[1][18][11] , \s_mux_signals[1][18][10] , 
        \s_mux_signals[1][18][9] , \s_mux_signals[1][18][8] , 
        \s_mux_signals[1][18][7] , \s_mux_signals[1][18][6] , 
        \s_mux_signals[1][18][5] , \s_mux_signals[1][18][4] , 
        \s_mux_signals[1][18][3] , \s_mux_signals[1][18][2] , 
        \s_mux_signals[1][18][1] , \s_mux_signals[1][18][0] }) );
  Mux_NBit_2x1_NBIT_IN32_111 MUX1_0_20 ( .port0({\s_mux_signals[0][20][31] , 
        \s_mux_signals[0][20][30] , \s_mux_signals[0][20][29] , 
        \s_mux_signals[0][20][28] , \s_mux_signals[0][20][27] , 
        \s_mux_signals[0][20][26] , \s_mux_signals[0][20][25] , 
        \s_mux_signals[0][20][24] , \s_mux_signals[0][20][23] , 
        \s_mux_signals[0][20][22] , \s_mux_signals[0][20][21] , 
        \s_mux_signals[0][20][20] , \s_mux_signals[0][20][19] , 
        \s_mux_signals[0][20][18] , \s_mux_signals[0][20][17] , 
        \s_mux_signals[0][20][16] , \s_mux_signals[0][20][15] , 
        \s_mux_signals[0][20][14] , \s_mux_signals[0][20][13] , 
        \s_mux_signals[0][20][12] , \s_mux_signals[0][20][11] , 
        \s_mux_signals[0][20][10] , \s_mux_signals[0][20][9] , 
        \s_mux_signals[0][20][8] , \s_mux_signals[0][20][7] , 
        \s_mux_signals[0][20][6] , \s_mux_signals[0][20][5] , 
        \s_mux_signals[0][20][4] , \s_mux_signals[0][20][3] , 
        \s_mux_signals[0][20][2] , \s_mux_signals[0][20][1] , 
        \s_mux_signals[0][20][0] }), .port1({\s_mux_signals[0][21][31] , 
        \s_mux_signals[0][21][30] , \s_mux_signals[0][21][29] , 
        \s_mux_signals[0][21][28] , \s_mux_signals[0][21][27] , 
        \s_mux_signals[0][21][26] , \s_mux_signals[0][21][25] , 
        \s_mux_signals[0][21][24] , \s_mux_signals[0][21][23] , 
        \s_mux_signals[0][21][22] , \s_mux_signals[0][21][21] , 
        \s_mux_signals[0][21][20] , \s_mux_signals[0][21][19] , 
        \s_mux_signals[0][21][18] , \s_mux_signals[0][21][17] , 
        \s_mux_signals[0][21][16] , \s_mux_signals[0][21][15] , 
        \s_mux_signals[0][21][14] , \s_mux_signals[0][21][13] , 
        \s_mux_signals[0][21][12] , \s_mux_signals[0][21][11] , 
        \s_mux_signals[0][21][10] , \s_mux_signals[0][21][9] , 
        \s_mux_signals[0][21][8] , \s_mux_signals[0][21][7] , 
        \s_mux_signals[0][21][6] , \s_mux_signals[0][21][5] , 
        \s_mux_signals[0][21][4] , \s_mux_signals[0][21][3] , 
        \s_mux_signals[0][21][2] , \s_mux_signals[0][21][1] , 
        \s_mux_signals[0][21][0] }), .sel(n12), .portY({
        \s_mux_signals[1][20][31] , \s_mux_signals[1][20][30] , 
        \s_mux_signals[1][20][29] , \s_mux_signals[1][20][28] , 
        \s_mux_signals[1][20][27] , \s_mux_signals[1][20][26] , 
        \s_mux_signals[1][20][25] , \s_mux_signals[1][20][24] , 
        \s_mux_signals[1][20][23] , \s_mux_signals[1][20][22] , 
        \s_mux_signals[1][20][21] , \s_mux_signals[1][20][20] , 
        \s_mux_signals[1][20][19] , \s_mux_signals[1][20][18] , 
        \s_mux_signals[1][20][17] , \s_mux_signals[1][20][16] , 
        \s_mux_signals[1][20][15] , \s_mux_signals[1][20][14] , 
        \s_mux_signals[1][20][13] , \s_mux_signals[1][20][12] , 
        \s_mux_signals[1][20][11] , \s_mux_signals[1][20][10] , 
        \s_mux_signals[1][20][9] , \s_mux_signals[1][20][8] , 
        \s_mux_signals[1][20][7] , \s_mux_signals[1][20][6] , 
        \s_mux_signals[1][20][5] , \s_mux_signals[1][20][4] , 
        \s_mux_signals[1][20][3] , \s_mux_signals[1][20][2] , 
        \s_mux_signals[1][20][1] , \s_mux_signals[1][20][0] }) );
  Mux_NBit_2x1_NBIT_IN32_110 MUX1_0_22 ( .port0({\s_mux_signals[0][22][31] , 
        \s_mux_signals[0][22][30] , \s_mux_signals[0][22][29] , 
        \s_mux_signals[0][22][28] , \s_mux_signals[0][22][27] , 
        \s_mux_signals[0][22][26] , \s_mux_signals[0][22][25] , 
        \s_mux_signals[0][22][24] , \s_mux_signals[0][22][23] , 
        \s_mux_signals[0][22][22] , \s_mux_signals[0][22][21] , 
        \s_mux_signals[0][22][20] , \s_mux_signals[0][22][19] , 
        \s_mux_signals[0][22][18] , \s_mux_signals[0][22][17] , 
        \s_mux_signals[0][22][16] , \s_mux_signals[0][22][15] , 
        \s_mux_signals[0][22][14] , \s_mux_signals[0][22][13] , 
        \s_mux_signals[0][22][12] , \s_mux_signals[0][22][11] , 
        \s_mux_signals[0][22][10] , \s_mux_signals[0][22][9] , 
        \s_mux_signals[0][22][8] , \s_mux_signals[0][22][7] , 
        \s_mux_signals[0][22][6] , \s_mux_signals[0][22][5] , 
        \s_mux_signals[0][22][4] , \s_mux_signals[0][22][3] , 
        \s_mux_signals[0][22][2] , \s_mux_signals[0][22][1] , 
        \s_mux_signals[0][22][0] }), .port1({\s_mux_signals[0][23][31] , 
        \s_mux_signals[0][23][30] , \s_mux_signals[0][23][29] , 
        \s_mux_signals[0][23][28] , \s_mux_signals[0][23][27] , 
        \s_mux_signals[0][23][26] , \s_mux_signals[0][23][25] , 
        \s_mux_signals[0][23][24] , \s_mux_signals[0][23][23] , 
        \s_mux_signals[0][23][22] , \s_mux_signals[0][23][21] , 
        \s_mux_signals[0][23][20] , \s_mux_signals[0][23][19] , 
        \s_mux_signals[0][23][18] , \s_mux_signals[0][23][17] , 
        \s_mux_signals[0][23][16] , \s_mux_signals[0][23][15] , 
        \s_mux_signals[0][23][14] , \s_mux_signals[0][23][13] , 
        \s_mux_signals[0][23][12] , \s_mux_signals[0][23][11] , 
        \s_mux_signals[0][23][10] , \s_mux_signals[0][23][9] , 
        \s_mux_signals[0][23][8] , \s_mux_signals[0][23][7] , 
        \s_mux_signals[0][23][6] , \s_mux_signals[0][23][5] , 
        \s_mux_signals[0][23][4] , \s_mux_signals[0][23][3] , 
        \s_mux_signals[0][23][2] , \s_mux_signals[0][23][1] , 
        \s_mux_signals[0][23][0] }), .sel(n12), .portY({
        \s_mux_signals[1][22][31] , \s_mux_signals[1][22][30] , 
        \s_mux_signals[1][22][29] , \s_mux_signals[1][22][28] , 
        \s_mux_signals[1][22][27] , \s_mux_signals[1][22][26] , 
        \s_mux_signals[1][22][25] , \s_mux_signals[1][22][24] , 
        \s_mux_signals[1][22][23] , \s_mux_signals[1][22][22] , 
        \s_mux_signals[1][22][21] , \s_mux_signals[1][22][20] , 
        \s_mux_signals[1][22][19] , \s_mux_signals[1][22][18] , 
        \s_mux_signals[1][22][17] , \s_mux_signals[1][22][16] , 
        \s_mux_signals[1][22][15] , \s_mux_signals[1][22][14] , 
        \s_mux_signals[1][22][13] , \s_mux_signals[1][22][12] , 
        \s_mux_signals[1][22][11] , \s_mux_signals[1][22][10] , 
        \s_mux_signals[1][22][9] , \s_mux_signals[1][22][8] , 
        \s_mux_signals[1][22][7] , \s_mux_signals[1][22][6] , 
        \s_mux_signals[1][22][5] , \s_mux_signals[1][22][4] , 
        \s_mux_signals[1][22][3] , \s_mux_signals[1][22][2] , 
        \s_mux_signals[1][22][1] , \s_mux_signals[1][22][0] }) );
  Mux_NBit_2x1_NBIT_IN32_109 MUX1_0_24 ( .port0({\s_mux_signals[0][24][31] , 
        \s_mux_signals[0][24][30] , \s_mux_signals[0][24][29] , 
        \s_mux_signals[0][24][28] , \s_mux_signals[0][24][27] , 
        \s_mux_signals[0][24][26] , \s_mux_signals[0][24][25] , 
        \s_mux_signals[0][24][24] , \s_mux_signals[0][24][23] , 
        \s_mux_signals[0][24][22] , \s_mux_signals[0][24][21] , 
        \s_mux_signals[0][24][20] , \s_mux_signals[0][24][19] , 
        \s_mux_signals[0][24][18] , \s_mux_signals[0][24][17] , 
        \s_mux_signals[0][24][16] , \s_mux_signals[0][24][15] , 
        \s_mux_signals[0][24][14] , \s_mux_signals[0][24][13] , 
        \s_mux_signals[0][24][12] , \s_mux_signals[0][24][11] , 
        \s_mux_signals[0][24][10] , \s_mux_signals[0][24][9] , 
        \s_mux_signals[0][24][8] , \s_mux_signals[0][24][7] , 
        \s_mux_signals[0][24][6] , \s_mux_signals[0][24][5] , 
        \s_mux_signals[0][24][4] , \s_mux_signals[0][24][3] , 
        \s_mux_signals[0][24][2] , \s_mux_signals[0][24][1] , 
        \s_mux_signals[0][24][0] }), .port1({\s_mux_signals[0][25][31] , 
        \s_mux_signals[0][25][30] , \s_mux_signals[0][25][29] , 
        \s_mux_signals[0][25][28] , \s_mux_signals[0][25][27] , 
        \s_mux_signals[0][25][26] , \s_mux_signals[0][25][25] , 
        \s_mux_signals[0][25][24] , \s_mux_signals[0][25][23] , 
        \s_mux_signals[0][25][22] , \s_mux_signals[0][25][21] , 
        \s_mux_signals[0][25][20] , \s_mux_signals[0][25][19] , 
        \s_mux_signals[0][25][18] , \s_mux_signals[0][25][17] , 
        \s_mux_signals[0][25][16] , \s_mux_signals[0][25][15] , 
        \s_mux_signals[0][25][14] , \s_mux_signals[0][25][13] , 
        \s_mux_signals[0][25][12] , \s_mux_signals[0][25][11] , 
        \s_mux_signals[0][25][10] , \s_mux_signals[0][25][9] , 
        \s_mux_signals[0][25][8] , \s_mux_signals[0][25][7] , 
        \s_mux_signals[0][25][6] , \s_mux_signals[0][25][5] , 
        \s_mux_signals[0][25][4] , \s_mux_signals[0][25][3] , 
        \s_mux_signals[0][25][2] , \s_mux_signals[0][25][1] , 
        \s_mux_signals[0][25][0] }), .sel(n12), .portY({
        \s_mux_signals[1][24][31] , \s_mux_signals[1][24][30] , 
        \s_mux_signals[1][24][29] , \s_mux_signals[1][24][28] , 
        \s_mux_signals[1][24][27] , \s_mux_signals[1][24][26] , 
        \s_mux_signals[1][24][25] , \s_mux_signals[1][24][24] , 
        \s_mux_signals[1][24][23] , \s_mux_signals[1][24][22] , 
        \s_mux_signals[1][24][21] , \s_mux_signals[1][24][20] , 
        \s_mux_signals[1][24][19] , \s_mux_signals[1][24][18] , 
        \s_mux_signals[1][24][17] , \s_mux_signals[1][24][16] , 
        \s_mux_signals[1][24][15] , \s_mux_signals[1][24][14] , 
        \s_mux_signals[1][24][13] , \s_mux_signals[1][24][12] , 
        \s_mux_signals[1][24][11] , \s_mux_signals[1][24][10] , 
        \s_mux_signals[1][24][9] , \s_mux_signals[1][24][8] , 
        \s_mux_signals[1][24][7] , \s_mux_signals[1][24][6] , 
        \s_mux_signals[1][24][5] , \s_mux_signals[1][24][4] , 
        \s_mux_signals[1][24][3] , \s_mux_signals[1][24][2] , 
        \s_mux_signals[1][24][1] , \s_mux_signals[1][24][0] }) );
  Mux_NBit_2x1_NBIT_IN32_108 MUX1_0_26 ( .port0({\s_mux_signals[0][26][31] , 
        \s_mux_signals[0][26][30] , \s_mux_signals[0][26][29] , 
        \s_mux_signals[0][26][28] , \s_mux_signals[0][26][27] , 
        \s_mux_signals[0][26][26] , \s_mux_signals[0][26][25] , 
        \s_mux_signals[0][26][24] , \s_mux_signals[0][26][23] , 
        \s_mux_signals[0][26][22] , \s_mux_signals[0][26][21] , 
        \s_mux_signals[0][26][20] , \s_mux_signals[0][26][19] , 
        \s_mux_signals[0][26][18] , \s_mux_signals[0][26][17] , 
        \s_mux_signals[0][26][16] , \s_mux_signals[0][26][15] , 
        \s_mux_signals[0][26][14] , \s_mux_signals[0][26][13] , 
        \s_mux_signals[0][26][12] , \s_mux_signals[0][26][11] , 
        \s_mux_signals[0][26][10] , \s_mux_signals[0][26][9] , 
        \s_mux_signals[0][26][8] , \s_mux_signals[0][26][7] , 
        \s_mux_signals[0][26][6] , \s_mux_signals[0][26][5] , 
        \s_mux_signals[0][26][4] , \s_mux_signals[0][26][3] , 
        \s_mux_signals[0][26][2] , \s_mux_signals[0][26][1] , 
        \s_mux_signals[0][26][0] }), .port1({\s_mux_signals[0][27][31] , 
        \s_mux_signals[0][27][30] , \s_mux_signals[0][27][29] , 
        \s_mux_signals[0][27][28] , \s_mux_signals[0][27][27] , 
        \s_mux_signals[0][27][26] , \s_mux_signals[0][27][25] , 
        \s_mux_signals[0][27][24] , \s_mux_signals[0][27][23] , 
        \s_mux_signals[0][27][22] , \s_mux_signals[0][27][21] , 
        \s_mux_signals[0][27][20] , \s_mux_signals[0][27][19] , 
        \s_mux_signals[0][27][18] , \s_mux_signals[0][27][17] , 
        \s_mux_signals[0][27][16] , \s_mux_signals[0][27][15] , 
        \s_mux_signals[0][27][14] , \s_mux_signals[0][27][13] , 
        \s_mux_signals[0][27][12] , \s_mux_signals[0][27][11] , 
        \s_mux_signals[0][27][10] , \s_mux_signals[0][27][9] , 
        \s_mux_signals[0][27][8] , \s_mux_signals[0][27][7] , 
        \s_mux_signals[0][27][6] , \s_mux_signals[0][27][5] , 
        \s_mux_signals[0][27][4] , \s_mux_signals[0][27][3] , 
        \s_mux_signals[0][27][2] , \s_mux_signals[0][27][1] , 
        \s_mux_signals[0][27][0] }), .sel(n12), .portY({
        \s_mux_signals[1][26][31] , \s_mux_signals[1][26][30] , 
        \s_mux_signals[1][26][29] , \s_mux_signals[1][26][28] , 
        \s_mux_signals[1][26][27] , \s_mux_signals[1][26][26] , 
        \s_mux_signals[1][26][25] , \s_mux_signals[1][26][24] , 
        \s_mux_signals[1][26][23] , \s_mux_signals[1][26][22] , 
        \s_mux_signals[1][26][21] , \s_mux_signals[1][26][20] , 
        \s_mux_signals[1][26][19] , \s_mux_signals[1][26][18] , 
        \s_mux_signals[1][26][17] , \s_mux_signals[1][26][16] , 
        \s_mux_signals[1][26][15] , \s_mux_signals[1][26][14] , 
        \s_mux_signals[1][26][13] , \s_mux_signals[1][26][12] , 
        \s_mux_signals[1][26][11] , \s_mux_signals[1][26][10] , 
        \s_mux_signals[1][26][9] , \s_mux_signals[1][26][8] , 
        \s_mux_signals[1][26][7] , \s_mux_signals[1][26][6] , 
        \s_mux_signals[1][26][5] , \s_mux_signals[1][26][4] , 
        \s_mux_signals[1][26][3] , \s_mux_signals[1][26][2] , 
        \s_mux_signals[1][26][1] , \s_mux_signals[1][26][0] }) );
  Mux_NBit_2x1_NBIT_IN32_107 MUX1_0_28 ( .port0({\s_mux_signals[0][28][31] , 
        \s_mux_signals[0][28][30] , \s_mux_signals[0][28][29] , 
        \s_mux_signals[0][28][28] , \s_mux_signals[0][28][27] , 
        \s_mux_signals[0][28][26] , \s_mux_signals[0][28][25] , 
        \s_mux_signals[0][28][24] , \s_mux_signals[0][28][23] , 
        \s_mux_signals[0][28][22] , \s_mux_signals[0][28][21] , 
        \s_mux_signals[0][28][20] , \s_mux_signals[0][28][19] , 
        \s_mux_signals[0][28][18] , \s_mux_signals[0][28][17] , 
        \s_mux_signals[0][28][16] , \s_mux_signals[0][28][15] , 
        \s_mux_signals[0][28][14] , \s_mux_signals[0][28][13] , 
        \s_mux_signals[0][28][12] , \s_mux_signals[0][28][11] , 
        \s_mux_signals[0][28][10] , \s_mux_signals[0][28][9] , 
        \s_mux_signals[0][28][8] , \s_mux_signals[0][28][7] , 
        \s_mux_signals[0][28][6] , \s_mux_signals[0][28][5] , 
        \s_mux_signals[0][28][4] , \s_mux_signals[0][28][3] , 
        \s_mux_signals[0][28][2] , \s_mux_signals[0][28][1] , 
        \s_mux_signals[0][28][0] }), .port1({\s_mux_signals[0][29][31] , 
        \s_mux_signals[0][29][30] , \s_mux_signals[0][29][29] , 
        \s_mux_signals[0][29][28] , \s_mux_signals[0][29][27] , 
        \s_mux_signals[0][29][26] , \s_mux_signals[0][29][25] , 
        \s_mux_signals[0][29][24] , \s_mux_signals[0][29][23] , 
        \s_mux_signals[0][29][22] , \s_mux_signals[0][29][21] , 
        \s_mux_signals[0][29][20] , \s_mux_signals[0][29][19] , 
        \s_mux_signals[0][29][18] , \s_mux_signals[0][29][17] , 
        \s_mux_signals[0][29][16] , \s_mux_signals[0][29][15] , 
        \s_mux_signals[0][29][14] , \s_mux_signals[0][29][13] , 
        \s_mux_signals[0][29][12] , \s_mux_signals[0][29][11] , 
        \s_mux_signals[0][29][10] , \s_mux_signals[0][29][9] , 
        \s_mux_signals[0][29][8] , \s_mux_signals[0][29][7] , 
        \s_mux_signals[0][29][6] , \s_mux_signals[0][29][5] , 
        \s_mux_signals[0][29][4] , \s_mux_signals[0][29][3] , 
        \s_mux_signals[0][29][2] , \s_mux_signals[0][29][1] , 
        \s_mux_signals[0][29][0] }), .sel(n12), .portY({
        \s_mux_signals[1][28][31] , \s_mux_signals[1][28][30] , 
        \s_mux_signals[1][28][29] , \s_mux_signals[1][28][28] , 
        \s_mux_signals[1][28][27] , \s_mux_signals[1][28][26] , 
        \s_mux_signals[1][28][25] , \s_mux_signals[1][28][24] , 
        \s_mux_signals[1][28][23] , \s_mux_signals[1][28][22] , 
        \s_mux_signals[1][28][21] , \s_mux_signals[1][28][20] , 
        \s_mux_signals[1][28][19] , \s_mux_signals[1][28][18] , 
        \s_mux_signals[1][28][17] , \s_mux_signals[1][28][16] , 
        \s_mux_signals[1][28][15] , \s_mux_signals[1][28][14] , 
        \s_mux_signals[1][28][13] , \s_mux_signals[1][28][12] , 
        \s_mux_signals[1][28][11] , \s_mux_signals[1][28][10] , 
        \s_mux_signals[1][28][9] , \s_mux_signals[1][28][8] , 
        \s_mux_signals[1][28][7] , \s_mux_signals[1][28][6] , 
        \s_mux_signals[1][28][5] , \s_mux_signals[1][28][4] , 
        \s_mux_signals[1][28][3] , \s_mux_signals[1][28][2] , 
        \s_mux_signals[1][28][1] , \s_mux_signals[1][28][0] }) );
  Mux_NBit_2x1_NBIT_IN32_106 MUX1_0_30 ( .port0({\s_mux_signals[0][30][31] , 
        \s_mux_signals[0][30][30] , \s_mux_signals[0][30][29] , 
        \s_mux_signals[0][30][28] , \s_mux_signals[0][30][27] , 
        \s_mux_signals[0][30][26] , \s_mux_signals[0][30][25] , 
        \s_mux_signals[0][30][24] , \s_mux_signals[0][30][23] , 
        \s_mux_signals[0][30][22] , \s_mux_signals[0][30][21] , 
        \s_mux_signals[0][30][20] , \s_mux_signals[0][30][19] , 
        \s_mux_signals[0][30][18] , \s_mux_signals[0][30][17] , 
        \s_mux_signals[0][30][16] , \s_mux_signals[0][30][15] , 
        \s_mux_signals[0][30][14] , \s_mux_signals[0][30][13] , 
        \s_mux_signals[0][30][12] , \s_mux_signals[0][30][11] , 
        \s_mux_signals[0][30][10] , \s_mux_signals[0][30][9] , 
        \s_mux_signals[0][30][8] , \s_mux_signals[0][30][7] , 
        \s_mux_signals[0][30][6] , \s_mux_signals[0][30][5] , 
        \s_mux_signals[0][30][4] , \s_mux_signals[0][30][3] , 
        \s_mux_signals[0][30][2] , \s_mux_signals[0][30][1] , 
        \s_mux_signals[0][30][0] }), .port1({\s_mux_signals[0][31][31] , 
        \s_mux_signals[0][31][30] , \s_mux_signals[0][31][29] , 
        \s_mux_signals[0][31][28] , \s_mux_signals[0][31][27] , 
        \s_mux_signals[0][31][26] , \s_mux_signals[0][31][25] , 
        \s_mux_signals[0][31][24] , \s_mux_signals[0][31][23] , 
        \s_mux_signals[0][31][22] , \s_mux_signals[0][31][21] , 
        \s_mux_signals[0][31][20] , \s_mux_signals[0][31][19] , 
        \s_mux_signals[0][31][18] , \s_mux_signals[0][31][17] , 
        \s_mux_signals[0][31][16] , \s_mux_signals[0][31][15] , 
        \s_mux_signals[0][31][14] , \s_mux_signals[0][31][13] , 
        \s_mux_signals[0][31][12] , \s_mux_signals[0][31][11] , 
        \s_mux_signals[0][31][10] , \s_mux_signals[0][31][9] , 
        \s_mux_signals[0][31][8] , \s_mux_signals[0][31][7] , 
        \s_mux_signals[0][31][6] , \s_mux_signals[0][31][5] , 
        \s_mux_signals[0][31][4] , \s_mux_signals[0][31][3] , 
        \s_mux_signals[0][31][2] , \s_mux_signals[0][31][1] , 
        \s_mux_signals[0][31][0] }), .sel(n13), .portY({
        \s_mux_signals[1][30][31] , \s_mux_signals[1][30][30] , 
        \s_mux_signals[1][30][29] , \s_mux_signals[1][30][28] , 
        \s_mux_signals[1][30][27] , \s_mux_signals[1][30][26] , 
        \s_mux_signals[1][30][25] , \s_mux_signals[1][30][24] , 
        \s_mux_signals[1][30][23] , \s_mux_signals[1][30][22] , 
        \s_mux_signals[1][30][21] , \s_mux_signals[1][30][20] , 
        \s_mux_signals[1][30][19] , \s_mux_signals[1][30][18] , 
        \s_mux_signals[1][30][17] , \s_mux_signals[1][30][16] , 
        \s_mux_signals[1][30][15] , \s_mux_signals[1][30][14] , 
        \s_mux_signals[1][30][13] , \s_mux_signals[1][30][12] , 
        \s_mux_signals[1][30][11] , \s_mux_signals[1][30][10] , 
        \s_mux_signals[1][30][9] , \s_mux_signals[1][30][8] , 
        \s_mux_signals[1][30][7] , \s_mux_signals[1][30][6] , 
        \s_mux_signals[1][30][5] , \s_mux_signals[1][30][4] , 
        \s_mux_signals[1][30][3] , \s_mux_signals[1][30][2] , 
        \s_mux_signals[1][30][1] , \s_mux_signals[1][30][0] }) );
  Mux_NBit_2x1_NBIT_IN32_105 MUX1_1_0 ( .port0({\s_mux_signals[1][0][31] , 
        \s_mux_signals[1][0][30] , \s_mux_signals[1][0][29] , 
        \s_mux_signals[1][0][28] , \s_mux_signals[1][0][27] , 
        \s_mux_signals[1][0][26] , \s_mux_signals[1][0][25] , 
        \s_mux_signals[1][0][24] , \s_mux_signals[1][0][23] , 
        \s_mux_signals[1][0][22] , \s_mux_signals[1][0][21] , 
        \s_mux_signals[1][0][20] , \s_mux_signals[1][0][19] , 
        \s_mux_signals[1][0][18] , \s_mux_signals[1][0][17] , 
        \s_mux_signals[1][0][16] , \s_mux_signals[1][0][15] , 
        \s_mux_signals[1][0][14] , \s_mux_signals[1][0][13] , 
        \s_mux_signals[1][0][12] , \s_mux_signals[1][0][11] , 
        \s_mux_signals[1][0][10] , \s_mux_signals[1][0][9] , 
        \s_mux_signals[1][0][8] , \s_mux_signals[1][0][7] , 
        \s_mux_signals[1][0][6] , \s_mux_signals[1][0][5] , 
        \s_mux_signals[1][0][4] , \s_mux_signals[1][0][3] , 
        \s_mux_signals[1][0][2] , \s_mux_signals[1][0][1] , 
        \s_mux_signals[1][0][0] }), .port1({\s_mux_signals[1][2][31] , 
        \s_mux_signals[1][2][30] , \s_mux_signals[1][2][29] , 
        \s_mux_signals[1][2][28] , \s_mux_signals[1][2][27] , 
        \s_mux_signals[1][2][26] , \s_mux_signals[1][2][25] , 
        \s_mux_signals[1][2][24] , \s_mux_signals[1][2][23] , 
        \s_mux_signals[1][2][22] , \s_mux_signals[1][2][21] , 
        \s_mux_signals[1][2][20] , \s_mux_signals[1][2][19] , 
        \s_mux_signals[1][2][18] , \s_mux_signals[1][2][17] , 
        \s_mux_signals[1][2][16] , \s_mux_signals[1][2][15] , 
        \s_mux_signals[1][2][14] , \s_mux_signals[1][2][13] , 
        \s_mux_signals[1][2][12] , \s_mux_signals[1][2][11] , 
        \s_mux_signals[1][2][10] , \s_mux_signals[1][2][9] , 
        \s_mux_signals[1][2][8] , \s_mux_signals[1][2][7] , 
        \s_mux_signals[1][2][6] , \s_mux_signals[1][2][5] , 
        \s_mux_signals[1][2][4] , \s_mux_signals[1][2][3] , 
        \s_mux_signals[1][2][2] , \s_mux_signals[1][2][1] , 
        \s_mux_signals[1][2][0] }), .sel(n23), .portY({
        \s_mux_signals[2][0][31] , \s_mux_signals[2][0][30] , 
        \s_mux_signals[2][0][29] , \s_mux_signals[2][0][28] , 
        \s_mux_signals[2][0][27] , \s_mux_signals[2][0][26] , 
        \s_mux_signals[2][0][25] , \s_mux_signals[2][0][24] , 
        \s_mux_signals[2][0][23] , \s_mux_signals[2][0][22] , 
        \s_mux_signals[2][0][21] , \s_mux_signals[2][0][20] , 
        \s_mux_signals[2][0][19] , \s_mux_signals[2][0][18] , 
        \s_mux_signals[2][0][17] , \s_mux_signals[2][0][16] , 
        \s_mux_signals[2][0][15] , \s_mux_signals[2][0][14] , 
        \s_mux_signals[2][0][13] , \s_mux_signals[2][0][12] , 
        \s_mux_signals[2][0][11] , \s_mux_signals[2][0][10] , 
        \s_mux_signals[2][0][9] , \s_mux_signals[2][0][8] , 
        \s_mux_signals[2][0][7] , \s_mux_signals[2][0][6] , 
        \s_mux_signals[2][0][5] , \s_mux_signals[2][0][4] , 
        \s_mux_signals[2][0][3] , \s_mux_signals[2][0][2] , 
        \s_mux_signals[2][0][1] , \s_mux_signals[2][0][0] }) );
  Mux_NBit_2x1_NBIT_IN32_104 MUX1_1_4 ( .port0({\s_mux_signals[1][4][31] , 
        \s_mux_signals[1][4][30] , \s_mux_signals[1][4][29] , 
        \s_mux_signals[1][4][28] , \s_mux_signals[1][4][27] , 
        \s_mux_signals[1][4][26] , \s_mux_signals[1][4][25] , 
        \s_mux_signals[1][4][24] , \s_mux_signals[1][4][23] , 
        \s_mux_signals[1][4][22] , \s_mux_signals[1][4][21] , 
        \s_mux_signals[1][4][20] , \s_mux_signals[1][4][19] , 
        \s_mux_signals[1][4][18] , \s_mux_signals[1][4][17] , 
        \s_mux_signals[1][4][16] , \s_mux_signals[1][4][15] , 
        \s_mux_signals[1][4][14] , \s_mux_signals[1][4][13] , 
        \s_mux_signals[1][4][12] , \s_mux_signals[1][4][11] , 
        \s_mux_signals[1][4][10] , \s_mux_signals[1][4][9] , 
        \s_mux_signals[1][4][8] , \s_mux_signals[1][4][7] , 
        \s_mux_signals[1][4][6] , \s_mux_signals[1][4][5] , 
        \s_mux_signals[1][4][4] , \s_mux_signals[1][4][3] , 
        \s_mux_signals[1][4][2] , \s_mux_signals[1][4][1] , 
        \s_mux_signals[1][4][0] }), .port1({\s_mux_signals[1][6][31] , 
        \s_mux_signals[1][6][30] , \s_mux_signals[1][6][29] , 
        \s_mux_signals[1][6][28] , \s_mux_signals[1][6][27] , 
        \s_mux_signals[1][6][26] , \s_mux_signals[1][6][25] , 
        \s_mux_signals[1][6][24] , \s_mux_signals[1][6][23] , 
        \s_mux_signals[1][6][22] , \s_mux_signals[1][6][21] , 
        \s_mux_signals[1][6][20] , \s_mux_signals[1][6][19] , 
        \s_mux_signals[1][6][18] , \s_mux_signals[1][6][17] , 
        \s_mux_signals[1][6][16] , \s_mux_signals[1][6][15] , 
        \s_mux_signals[1][6][14] , \s_mux_signals[1][6][13] , 
        \s_mux_signals[1][6][12] , \s_mux_signals[1][6][11] , 
        \s_mux_signals[1][6][10] , \s_mux_signals[1][6][9] , 
        \s_mux_signals[1][6][8] , \s_mux_signals[1][6][7] , 
        \s_mux_signals[1][6][6] , \s_mux_signals[1][6][5] , 
        \s_mux_signals[1][6][4] , \s_mux_signals[1][6][3] , 
        \s_mux_signals[1][6][2] , \s_mux_signals[1][6][1] , 
        \s_mux_signals[1][6][0] }), .sel(n23), .portY({
        \s_mux_signals[2][4][31] , \s_mux_signals[2][4][30] , 
        \s_mux_signals[2][4][29] , \s_mux_signals[2][4][28] , 
        \s_mux_signals[2][4][27] , \s_mux_signals[2][4][26] , 
        \s_mux_signals[2][4][25] , \s_mux_signals[2][4][24] , 
        \s_mux_signals[2][4][23] , \s_mux_signals[2][4][22] , 
        \s_mux_signals[2][4][21] , \s_mux_signals[2][4][20] , 
        \s_mux_signals[2][4][19] , \s_mux_signals[2][4][18] , 
        \s_mux_signals[2][4][17] , \s_mux_signals[2][4][16] , 
        \s_mux_signals[2][4][15] , \s_mux_signals[2][4][14] , 
        \s_mux_signals[2][4][13] , \s_mux_signals[2][4][12] , 
        \s_mux_signals[2][4][11] , \s_mux_signals[2][4][10] , 
        \s_mux_signals[2][4][9] , \s_mux_signals[2][4][8] , 
        \s_mux_signals[2][4][7] , \s_mux_signals[2][4][6] , 
        \s_mux_signals[2][4][5] , \s_mux_signals[2][4][4] , 
        \s_mux_signals[2][4][3] , \s_mux_signals[2][4][2] , 
        \s_mux_signals[2][4][1] , \s_mux_signals[2][4][0] }) );
  Mux_NBit_2x1_NBIT_IN32_103 MUX1_1_8 ( .port0({\s_mux_signals[1][8][31] , 
        \s_mux_signals[1][8][30] , \s_mux_signals[1][8][29] , 
        \s_mux_signals[1][8][28] , \s_mux_signals[1][8][27] , 
        \s_mux_signals[1][8][26] , \s_mux_signals[1][8][25] , 
        \s_mux_signals[1][8][24] , \s_mux_signals[1][8][23] , 
        \s_mux_signals[1][8][22] , \s_mux_signals[1][8][21] , 
        \s_mux_signals[1][8][20] , \s_mux_signals[1][8][19] , 
        \s_mux_signals[1][8][18] , \s_mux_signals[1][8][17] , 
        \s_mux_signals[1][8][16] , \s_mux_signals[1][8][15] , 
        \s_mux_signals[1][8][14] , \s_mux_signals[1][8][13] , 
        \s_mux_signals[1][8][12] , \s_mux_signals[1][8][11] , 
        \s_mux_signals[1][8][10] , \s_mux_signals[1][8][9] , 
        \s_mux_signals[1][8][8] , \s_mux_signals[1][8][7] , 
        \s_mux_signals[1][8][6] , \s_mux_signals[1][8][5] , 
        \s_mux_signals[1][8][4] , \s_mux_signals[1][8][3] , 
        \s_mux_signals[1][8][2] , \s_mux_signals[1][8][1] , 
        \s_mux_signals[1][8][0] }), .port1({\s_mux_signals[1][10][31] , 
        \s_mux_signals[1][10][30] , \s_mux_signals[1][10][29] , 
        \s_mux_signals[1][10][28] , \s_mux_signals[1][10][27] , 
        \s_mux_signals[1][10][26] , \s_mux_signals[1][10][25] , 
        \s_mux_signals[1][10][24] , \s_mux_signals[1][10][23] , 
        \s_mux_signals[1][10][22] , \s_mux_signals[1][10][21] , 
        \s_mux_signals[1][10][20] , \s_mux_signals[1][10][19] , 
        \s_mux_signals[1][10][18] , \s_mux_signals[1][10][17] , 
        \s_mux_signals[1][10][16] , \s_mux_signals[1][10][15] , 
        \s_mux_signals[1][10][14] , \s_mux_signals[1][10][13] , 
        \s_mux_signals[1][10][12] , \s_mux_signals[1][10][11] , 
        \s_mux_signals[1][10][10] , \s_mux_signals[1][10][9] , 
        \s_mux_signals[1][10][8] , \s_mux_signals[1][10][7] , 
        \s_mux_signals[1][10][6] , \s_mux_signals[1][10][5] , 
        \s_mux_signals[1][10][4] , \s_mux_signals[1][10][3] , 
        \s_mux_signals[1][10][2] , \s_mux_signals[1][10][1] , 
        \s_mux_signals[1][10][0] }), .sel(n23), .portY({
        \s_mux_signals[2][8][31] , \s_mux_signals[2][8][30] , 
        \s_mux_signals[2][8][29] , \s_mux_signals[2][8][28] , 
        \s_mux_signals[2][8][27] , \s_mux_signals[2][8][26] , 
        \s_mux_signals[2][8][25] , \s_mux_signals[2][8][24] , 
        \s_mux_signals[2][8][23] , \s_mux_signals[2][8][22] , 
        \s_mux_signals[2][8][21] , \s_mux_signals[2][8][20] , 
        \s_mux_signals[2][8][19] , \s_mux_signals[2][8][18] , 
        \s_mux_signals[2][8][17] , \s_mux_signals[2][8][16] , 
        \s_mux_signals[2][8][15] , \s_mux_signals[2][8][14] , 
        \s_mux_signals[2][8][13] , \s_mux_signals[2][8][12] , 
        \s_mux_signals[2][8][11] , \s_mux_signals[2][8][10] , 
        \s_mux_signals[2][8][9] , \s_mux_signals[2][8][8] , 
        \s_mux_signals[2][8][7] , \s_mux_signals[2][8][6] , 
        \s_mux_signals[2][8][5] , \s_mux_signals[2][8][4] , 
        \s_mux_signals[2][8][3] , \s_mux_signals[2][8][2] , 
        \s_mux_signals[2][8][1] , \s_mux_signals[2][8][0] }) );
  Mux_NBit_2x1_NBIT_IN32_102 MUX1_1_12 ( .port0({\s_mux_signals[1][12][31] , 
        \s_mux_signals[1][12][30] , \s_mux_signals[1][12][29] , 
        \s_mux_signals[1][12][28] , \s_mux_signals[1][12][27] , 
        \s_mux_signals[1][12][26] , \s_mux_signals[1][12][25] , 
        \s_mux_signals[1][12][24] , \s_mux_signals[1][12][23] , 
        \s_mux_signals[1][12][22] , \s_mux_signals[1][12][21] , 
        \s_mux_signals[1][12][20] , \s_mux_signals[1][12][19] , 
        \s_mux_signals[1][12][18] , \s_mux_signals[1][12][17] , 
        \s_mux_signals[1][12][16] , \s_mux_signals[1][12][15] , 
        \s_mux_signals[1][12][14] , \s_mux_signals[1][12][13] , 
        \s_mux_signals[1][12][12] , \s_mux_signals[1][12][11] , 
        \s_mux_signals[1][12][10] , \s_mux_signals[1][12][9] , 
        \s_mux_signals[1][12][8] , \s_mux_signals[1][12][7] , 
        \s_mux_signals[1][12][6] , \s_mux_signals[1][12][5] , 
        \s_mux_signals[1][12][4] , \s_mux_signals[1][12][3] , 
        \s_mux_signals[1][12][2] , \s_mux_signals[1][12][1] , 
        \s_mux_signals[1][12][0] }), .port1({\s_mux_signals[1][14][31] , 
        \s_mux_signals[1][14][30] , \s_mux_signals[1][14][29] , 
        \s_mux_signals[1][14][28] , \s_mux_signals[1][14][27] , 
        \s_mux_signals[1][14][26] , \s_mux_signals[1][14][25] , 
        \s_mux_signals[1][14][24] , \s_mux_signals[1][14][23] , 
        \s_mux_signals[1][14][22] , \s_mux_signals[1][14][21] , 
        \s_mux_signals[1][14][20] , \s_mux_signals[1][14][19] , 
        \s_mux_signals[1][14][18] , \s_mux_signals[1][14][17] , 
        \s_mux_signals[1][14][16] , \s_mux_signals[1][14][15] , 
        \s_mux_signals[1][14][14] , \s_mux_signals[1][14][13] , 
        \s_mux_signals[1][14][12] , \s_mux_signals[1][14][11] , 
        \s_mux_signals[1][14][10] , \s_mux_signals[1][14][9] , 
        \s_mux_signals[1][14][8] , \s_mux_signals[1][14][7] , 
        \s_mux_signals[1][14][6] , \s_mux_signals[1][14][5] , 
        \s_mux_signals[1][14][4] , \s_mux_signals[1][14][3] , 
        \s_mux_signals[1][14][2] , \s_mux_signals[1][14][1] , 
        \s_mux_signals[1][14][0] }), .sel(n24), .portY({
        \s_mux_signals[2][12][31] , \s_mux_signals[2][12][30] , 
        \s_mux_signals[2][12][29] , \s_mux_signals[2][12][28] , 
        \s_mux_signals[2][12][27] , \s_mux_signals[2][12][26] , 
        \s_mux_signals[2][12][25] , \s_mux_signals[2][12][24] , 
        \s_mux_signals[2][12][23] , \s_mux_signals[2][12][22] , 
        \s_mux_signals[2][12][21] , \s_mux_signals[2][12][20] , 
        \s_mux_signals[2][12][19] , \s_mux_signals[2][12][18] , 
        \s_mux_signals[2][12][17] , \s_mux_signals[2][12][16] , 
        \s_mux_signals[2][12][15] , \s_mux_signals[2][12][14] , 
        \s_mux_signals[2][12][13] , \s_mux_signals[2][12][12] , 
        \s_mux_signals[2][12][11] , \s_mux_signals[2][12][10] , 
        \s_mux_signals[2][12][9] , \s_mux_signals[2][12][8] , 
        \s_mux_signals[2][12][7] , \s_mux_signals[2][12][6] , 
        \s_mux_signals[2][12][5] , \s_mux_signals[2][12][4] , 
        \s_mux_signals[2][12][3] , \s_mux_signals[2][12][2] , 
        \s_mux_signals[2][12][1] , \s_mux_signals[2][12][0] }) );
  Mux_NBit_2x1_NBIT_IN32_101 MUX1_1_16 ( .port0({\s_mux_signals[1][16][31] , 
        \s_mux_signals[1][16][30] , \s_mux_signals[1][16][29] , 
        \s_mux_signals[1][16][28] , \s_mux_signals[1][16][27] , 
        \s_mux_signals[1][16][26] , \s_mux_signals[1][16][25] , 
        \s_mux_signals[1][16][24] , \s_mux_signals[1][16][23] , 
        \s_mux_signals[1][16][22] , \s_mux_signals[1][16][21] , 
        \s_mux_signals[1][16][20] , \s_mux_signals[1][16][19] , 
        \s_mux_signals[1][16][18] , \s_mux_signals[1][16][17] , 
        \s_mux_signals[1][16][16] , \s_mux_signals[1][16][15] , 
        \s_mux_signals[1][16][14] , \s_mux_signals[1][16][13] , 
        \s_mux_signals[1][16][12] , \s_mux_signals[1][16][11] , 
        \s_mux_signals[1][16][10] , \s_mux_signals[1][16][9] , 
        \s_mux_signals[1][16][8] , \s_mux_signals[1][16][7] , 
        \s_mux_signals[1][16][6] , \s_mux_signals[1][16][5] , 
        \s_mux_signals[1][16][4] , \s_mux_signals[1][16][3] , 
        \s_mux_signals[1][16][2] , \s_mux_signals[1][16][1] , 
        \s_mux_signals[1][16][0] }), .port1({\s_mux_signals[1][18][31] , 
        \s_mux_signals[1][18][30] , \s_mux_signals[1][18][29] , 
        \s_mux_signals[1][18][28] , \s_mux_signals[1][18][27] , 
        \s_mux_signals[1][18][26] , \s_mux_signals[1][18][25] , 
        \s_mux_signals[1][18][24] , \s_mux_signals[1][18][23] , 
        \s_mux_signals[1][18][22] , \s_mux_signals[1][18][21] , 
        \s_mux_signals[1][18][20] , \s_mux_signals[1][18][19] , 
        \s_mux_signals[1][18][18] , \s_mux_signals[1][18][17] , 
        \s_mux_signals[1][18][16] , \s_mux_signals[1][18][15] , 
        \s_mux_signals[1][18][14] , \s_mux_signals[1][18][13] , 
        \s_mux_signals[1][18][12] , \s_mux_signals[1][18][11] , 
        \s_mux_signals[1][18][10] , \s_mux_signals[1][18][9] , 
        \s_mux_signals[1][18][8] , \s_mux_signals[1][18][7] , 
        \s_mux_signals[1][18][6] , \s_mux_signals[1][18][5] , 
        \s_mux_signals[1][18][4] , \s_mux_signals[1][18][3] , 
        \s_mux_signals[1][18][2] , \s_mux_signals[1][18][1] , 
        \s_mux_signals[1][18][0] }), .sel(n24), .portY({
        \s_mux_signals[2][16][31] , \s_mux_signals[2][16][30] , 
        \s_mux_signals[2][16][29] , \s_mux_signals[2][16][28] , 
        \s_mux_signals[2][16][27] , \s_mux_signals[2][16][26] , 
        \s_mux_signals[2][16][25] , \s_mux_signals[2][16][24] , 
        \s_mux_signals[2][16][23] , \s_mux_signals[2][16][22] , 
        \s_mux_signals[2][16][21] , \s_mux_signals[2][16][20] , 
        \s_mux_signals[2][16][19] , \s_mux_signals[2][16][18] , 
        \s_mux_signals[2][16][17] , \s_mux_signals[2][16][16] , 
        \s_mux_signals[2][16][15] , \s_mux_signals[2][16][14] , 
        \s_mux_signals[2][16][13] , \s_mux_signals[2][16][12] , 
        \s_mux_signals[2][16][11] , \s_mux_signals[2][16][10] , 
        \s_mux_signals[2][16][9] , \s_mux_signals[2][16][8] , 
        \s_mux_signals[2][16][7] , \s_mux_signals[2][16][6] , 
        \s_mux_signals[2][16][5] , \s_mux_signals[2][16][4] , 
        \s_mux_signals[2][16][3] , \s_mux_signals[2][16][2] , 
        \s_mux_signals[2][16][1] , \s_mux_signals[2][16][0] }) );
  Mux_NBit_2x1_NBIT_IN32_100 MUX1_1_20 ( .port0({\s_mux_signals[1][20][31] , 
        \s_mux_signals[1][20][30] , \s_mux_signals[1][20][29] , 
        \s_mux_signals[1][20][28] , \s_mux_signals[1][20][27] , 
        \s_mux_signals[1][20][26] , \s_mux_signals[1][20][25] , 
        \s_mux_signals[1][20][24] , \s_mux_signals[1][20][23] , 
        \s_mux_signals[1][20][22] , \s_mux_signals[1][20][21] , 
        \s_mux_signals[1][20][20] , \s_mux_signals[1][20][19] , 
        \s_mux_signals[1][20][18] , \s_mux_signals[1][20][17] , 
        \s_mux_signals[1][20][16] , \s_mux_signals[1][20][15] , 
        \s_mux_signals[1][20][14] , \s_mux_signals[1][20][13] , 
        \s_mux_signals[1][20][12] , \s_mux_signals[1][20][11] , 
        \s_mux_signals[1][20][10] , \s_mux_signals[1][20][9] , 
        \s_mux_signals[1][20][8] , \s_mux_signals[1][20][7] , 
        \s_mux_signals[1][20][6] , \s_mux_signals[1][20][5] , 
        \s_mux_signals[1][20][4] , \s_mux_signals[1][20][3] , 
        \s_mux_signals[1][20][2] , \s_mux_signals[1][20][1] , 
        \s_mux_signals[1][20][0] }), .port1({\s_mux_signals[1][22][31] , 
        \s_mux_signals[1][22][30] , \s_mux_signals[1][22][29] , 
        \s_mux_signals[1][22][28] , \s_mux_signals[1][22][27] , 
        \s_mux_signals[1][22][26] , \s_mux_signals[1][22][25] , 
        \s_mux_signals[1][22][24] , \s_mux_signals[1][22][23] , 
        \s_mux_signals[1][22][22] , \s_mux_signals[1][22][21] , 
        \s_mux_signals[1][22][20] , \s_mux_signals[1][22][19] , 
        \s_mux_signals[1][22][18] , \s_mux_signals[1][22][17] , 
        \s_mux_signals[1][22][16] , \s_mux_signals[1][22][15] , 
        \s_mux_signals[1][22][14] , \s_mux_signals[1][22][13] , 
        \s_mux_signals[1][22][12] , \s_mux_signals[1][22][11] , 
        \s_mux_signals[1][22][10] , \s_mux_signals[1][22][9] , 
        \s_mux_signals[1][22][8] , \s_mux_signals[1][22][7] , 
        \s_mux_signals[1][22][6] , \s_mux_signals[1][22][5] , 
        \s_mux_signals[1][22][4] , \s_mux_signals[1][22][3] , 
        \s_mux_signals[1][22][2] , \s_mux_signals[1][22][1] , 
        \s_mux_signals[1][22][0] }), .sel(n24), .portY({
        \s_mux_signals[2][20][31] , \s_mux_signals[2][20][30] , 
        \s_mux_signals[2][20][29] , \s_mux_signals[2][20][28] , 
        \s_mux_signals[2][20][27] , \s_mux_signals[2][20][26] , 
        \s_mux_signals[2][20][25] , \s_mux_signals[2][20][24] , 
        \s_mux_signals[2][20][23] , \s_mux_signals[2][20][22] , 
        \s_mux_signals[2][20][21] , \s_mux_signals[2][20][20] , 
        \s_mux_signals[2][20][19] , \s_mux_signals[2][20][18] , 
        \s_mux_signals[2][20][17] , \s_mux_signals[2][20][16] , 
        \s_mux_signals[2][20][15] , \s_mux_signals[2][20][14] , 
        \s_mux_signals[2][20][13] , \s_mux_signals[2][20][12] , 
        \s_mux_signals[2][20][11] , \s_mux_signals[2][20][10] , 
        \s_mux_signals[2][20][9] , \s_mux_signals[2][20][8] , 
        \s_mux_signals[2][20][7] , \s_mux_signals[2][20][6] , 
        \s_mux_signals[2][20][5] , \s_mux_signals[2][20][4] , 
        \s_mux_signals[2][20][3] , \s_mux_signals[2][20][2] , 
        \s_mux_signals[2][20][1] , \s_mux_signals[2][20][0] }) );
  Mux_NBit_2x1_NBIT_IN32_99 MUX1_1_24 ( .port0({\s_mux_signals[1][24][31] , 
        \s_mux_signals[1][24][30] , \s_mux_signals[1][24][29] , 
        \s_mux_signals[1][24][28] , \s_mux_signals[1][24][27] , 
        \s_mux_signals[1][24][26] , \s_mux_signals[1][24][25] , 
        \s_mux_signals[1][24][24] , \s_mux_signals[1][24][23] , 
        \s_mux_signals[1][24][22] , \s_mux_signals[1][24][21] , 
        \s_mux_signals[1][24][20] , \s_mux_signals[1][24][19] , 
        \s_mux_signals[1][24][18] , \s_mux_signals[1][24][17] , 
        \s_mux_signals[1][24][16] , \s_mux_signals[1][24][15] , 
        \s_mux_signals[1][24][14] , \s_mux_signals[1][24][13] , 
        \s_mux_signals[1][24][12] , \s_mux_signals[1][24][11] , 
        \s_mux_signals[1][24][10] , \s_mux_signals[1][24][9] , 
        \s_mux_signals[1][24][8] , \s_mux_signals[1][24][7] , 
        \s_mux_signals[1][24][6] , \s_mux_signals[1][24][5] , 
        \s_mux_signals[1][24][4] , \s_mux_signals[1][24][3] , 
        \s_mux_signals[1][24][2] , \s_mux_signals[1][24][1] , 
        \s_mux_signals[1][24][0] }), .port1({\s_mux_signals[1][26][31] , 
        \s_mux_signals[1][26][30] , \s_mux_signals[1][26][29] , 
        \s_mux_signals[1][26][28] , \s_mux_signals[1][26][27] , 
        \s_mux_signals[1][26][26] , \s_mux_signals[1][26][25] , 
        \s_mux_signals[1][26][24] , \s_mux_signals[1][26][23] , 
        \s_mux_signals[1][26][22] , \s_mux_signals[1][26][21] , 
        \s_mux_signals[1][26][20] , \s_mux_signals[1][26][19] , 
        \s_mux_signals[1][26][18] , \s_mux_signals[1][26][17] , 
        \s_mux_signals[1][26][16] , \s_mux_signals[1][26][15] , 
        \s_mux_signals[1][26][14] , \s_mux_signals[1][26][13] , 
        \s_mux_signals[1][26][12] , \s_mux_signals[1][26][11] , 
        \s_mux_signals[1][26][10] , \s_mux_signals[1][26][9] , 
        \s_mux_signals[1][26][8] , \s_mux_signals[1][26][7] , 
        \s_mux_signals[1][26][6] , \s_mux_signals[1][26][5] , 
        \s_mux_signals[1][26][4] , \s_mux_signals[1][26][3] , 
        \s_mux_signals[1][26][2] , \s_mux_signals[1][26][1] , 
        \s_mux_signals[1][26][0] }), .sel(n25), .portY({
        \s_mux_signals[2][24][31] , \s_mux_signals[2][24][30] , 
        \s_mux_signals[2][24][29] , \s_mux_signals[2][24][28] , 
        \s_mux_signals[2][24][27] , \s_mux_signals[2][24][26] , 
        \s_mux_signals[2][24][25] , \s_mux_signals[2][24][24] , 
        \s_mux_signals[2][24][23] , \s_mux_signals[2][24][22] , 
        \s_mux_signals[2][24][21] , \s_mux_signals[2][24][20] , 
        \s_mux_signals[2][24][19] , \s_mux_signals[2][24][18] , 
        \s_mux_signals[2][24][17] , \s_mux_signals[2][24][16] , 
        \s_mux_signals[2][24][15] , \s_mux_signals[2][24][14] , 
        \s_mux_signals[2][24][13] , \s_mux_signals[2][24][12] , 
        \s_mux_signals[2][24][11] , \s_mux_signals[2][24][10] , 
        \s_mux_signals[2][24][9] , \s_mux_signals[2][24][8] , 
        \s_mux_signals[2][24][7] , \s_mux_signals[2][24][6] , 
        \s_mux_signals[2][24][5] , \s_mux_signals[2][24][4] , 
        \s_mux_signals[2][24][3] , \s_mux_signals[2][24][2] , 
        \s_mux_signals[2][24][1] , \s_mux_signals[2][24][0] }) );
  Mux_NBit_2x1_NBIT_IN32_98 MUX1_1_28 ( .port0({\s_mux_signals[1][28][31] , 
        \s_mux_signals[1][28][30] , \s_mux_signals[1][28][29] , 
        \s_mux_signals[1][28][28] , \s_mux_signals[1][28][27] , 
        \s_mux_signals[1][28][26] , \s_mux_signals[1][28][25] , 
        \s_mux_signals[1][28][24] , \s_mux_signals[1][28][23] , 
        \s_mux_signals[1][28][22] , \s_mux_signals[1][28][21] , 
        \s_mux_signals[1][28][20] , \s_mux_signals[1][28][19] , 
        \s_mux_signals[1][28][18] , \s_mux_signals[1][28][17] , 
        \s_mux_signals[1][28][16] , \s_mux_signals[1][28][15] , 
        \s_mux_signals[1][28][14] , \s_mux_signals[1][28][13] , 
        \s_mux_signals[1][28][12] , \s_mux_signals[1][28][11] , 
        \s_mux_signals[1][28][10] , \s_mux_signals[1][28][9] , 
        \s_mux_signals[1][28][8] , \s_mux_signals[1][28][7] , 
        \s_mux_signals[1][28][6] , \s_mux_signals[1][28][5] , 
        \s_mux_signals[1][28][4] , \s_mux_signals[1][28][3] , 
        \s_mux_signals[1][28][2] , \s_mux_signals[1][28][1] , 
        \s_mux_signals[1][28][0] }), .port1({\s_mux_signals[1][30][31] , 
        \s_mux_signals[1][30][30] , \s_mux_signals[1][30][29] , 
        \s_mux_signals[1][30][28] , \s_mux_signals[1][30][27] , 
        \s_mux_signals[1][30][26] , \s_mux_signals[1][30][25] , 
        \s_mux_signals[1][30][24] , \s_mux_signals[1][30][23] , 
        \s_mux_signals[1][30][22] , \s_mux_signals[1][30][21] , 
        \s_mux_signals[1][30][20] , \s_mux_signals[1][30][19] , 
        \s_mux_signals[1][30][18] , \s_mux_signals[1][30][17] , 
        \s_mux_signals[1][30][16] , \s_mux_signals[1][30][15] , 
        \s_mux_signals[1][30][14] , \s_mux_signals[1][30][13] , 
        \s_mux_signals[1][30][12] , \s_mux_signals[1][30][11] , 
        \s_mux_signals[1][30][10] , \s_mux_signals[1][30][9] , 
        \s_mux_signals[1][30][8] , \s_mux_signals[1][30][7] , 
        \s_mux_signals[1][30][6] , \s_mux_signals[1][30][5] , 
        \s_mux_signals[1][30][4] , \s_mux_signals[1][30][3] , 
        \s_mux_signals[1][30][2] , \s_mux_signals[1][30][1] , 
        \s_mux_signals[1][30][0] }), .sel(n25), .portY({
        \s_mux_signals[2][28][31] , \s_mux_signals[2][28][30] , 
        \s_mux_signals[2][28][29] , \s_mux_signals[2][28][28] , 
        \s_mux_signals[2][28][27] , \s_mux_signals[2][28][26] , 
        \s_mux_signals[2][28][25] , \s_mux_signals[2][28][24] , 
        \s_mux_signals[2][28][23] , \s_mux_signals[2][28][22] , 
        \s_mux_signals[2][28][21] , \s_mux_signals[2][28][20] , 
        \s_mux_signals[2][28][19] , \s_mux_signals[2][28][18] , 
        \s_mux_signals[2][28][17] , \s_mux_signals[2][28][16] , 
        \s_mux_signals[2][28][15] , \s_mux_signals[2][28][14] , 
        \s_mux_signals[2][28][13] , \s_mux_signals[2][28][12] , 
        \s_mux_signals[2][28][11] , \s_mux_signals[2][28][10] , 
        \s_mux_signals[2][28][9] , \s_mux_signals[2][28][8] , 
        \s_mux_signals[2][28][7] , \s_mux_signals[2][28][6] , 
        \s_mux_signals[2][28][5] , \s_mux_signals[2][28][4] , 
        \s_mux_signals[2][28][3] , \s_mux_signals[2][28][2] , 
        \s_mux_signals[2][28][1] , \s_mux_signals[2][28][0] }) );
  Mux_NBit_2x1_NBIT_IN32_97 MUX1_2_0 ( .port0({\s_mux_signals[2][0][31] , 
        \s_mux_signals[2][0][30] , \s_mux_signals[2][0][29] , 
        \s_mux_signals[2][0][28] , \s_mux_signals[2][0][27] , 
        \s_mux_signals[2][0][26] , \s_mux_signals[2][0][25] , 
        \s_mux_signals[2][0][24] , \s_mux_signals[2][0][23] , 
        \s_mux_signals[2][0][22] , \s_mux_signals[2][0][21] , 
        \s_mux_signals[2][0][20] , \s_mux_signals[2][0][19] , 
        \s_mux_signals[2][0][18] , \s_mux_signals[2][0][17] , 
        \s_mux_signals[2][0][16] , \s_mux_signals[2][0][15] , 
        \s_mux_signals[2][0][14] , \s_mux_signals[2][0][13] , 
        \s_mux_signals[2][0][12] , \s_mux_signals[2][0][11] , 
        \s_mux_signals[2][0][10] , \s_mux_signals[2][0][9] , 
        \s_mux_signals[2][0][8] , \s_mux_signals[2][0][7] , 
        \s_mux_signals[2][0][6] , \s_mux_signals[2][0][5] , 
        \s_mux_signals[2][0][4] , \s_mux_signals[2][0][3] , 
        \s_mux_signals[2][0][2] , \s_mux_signals[2][0][1] , 
        \s_mux_signals[2][0][0] }), .port1({\s_mux_signals[2][4][31] , 
        \s_mux_signals[2][4][30] , \s_mux_signals[2][4][29] , 
        \s_mux_signals[2][4][28] , \s_mux_signals[2][4][27] , 
        \s_mux_signals[2][4][26] , \s_mux_signals[2][4][25] , 
        \s_mux_signals[2][4][24] , \s_mux_signals[2][4][23] , 
        \s_mux_signals[2][4][22] , \s_mux_signals[2][4][21] , 
        \s_mux_signals[2][4][20] , \s_mux_signals[2][4][19] , 
        \s_mux_signals[2][4][18] , \s_mux_signals[2][4][17] , 
        \s_mux_signals[2][4][16] , \s_mux_signals[2][4][15] , 
        \s_mux_signals[2][4][14] , \s_mux_signals[2][4][13] , 
        \s_mux_signals[2][4][12] , \s_mux_signals[2][4][11] , 
        \s_mux_signals[2][4][10] , \s_mux_signals[2][4][9] , 
        \s_mux_signals[2][4][8] , \s_mux_signals[2][4][7] , 
        \s_mux_signals[2][4][6] , \s_mux_signals[2][4][5] , 
        \s_mux_signals[2][4][4] , \s_mux_signals[2][4][3] , 
        \s_mux_signals[2][4][2] , \s_mux_signals[2][4][1] , 
        \s_mux_signals[2][4][0] }), .sel(n26), .portY({
        \s_mux_signals[3][0][31] , \s_mux_signals[3][0][30] , 
        \s_mux_signals[3][0][29] , \s_mux_signals[3][0][28] , 
        \s_mux_signals[3][0][27] , \s_mux_signals[3][0][26] , 
        \s_mux_signals[3][0][25] , \s_mux_signals[3][0][24] , 
        \s_mux_signals[3][0][23] , \s_mux_signals[3][0][22] , 
        \s_mux_signals[3][0][21] , \s_mux_signals[3][0][20] , 
        \s_mux_signals[3][0][19] , \s_mux_signals[3][0][18] , 
        \s_mux_signals[3][0][17] , \s_mux_signals[3][0][16] , 
        \s_mux_signals[3][0][15] , \s_mux_signals[3][0][14] , 
        \s_mux_signals[3][0][13] , \s_mux_signals[3][0][12] , 
        \s_mux_signals[3][0][11] , \s_mux_signals[3][0][10] , 
        \s_mux_signals[3][0][9] , \s_mux_signals[3][0][8] , 
        \s_mux_signals[3][0][7] , \s_mux_signals[3][0][6] , 
        \s_mux_signals[3][0][5] , \s_mux_signals[3][0][4] , 
        \s_mux_signals[3][0][3] , \s_mux_signals[3][0][2] , 
        \s_mux_signals[3][0][1] , \s_mux_signals[3][0][0] }) );
  Mux_NBit_2x1_NBIT_IN32_96 MUX1_2_8 ( .port0({\s_mux_signals[2][8][31] , 
        \s_mux_signals[2][8][30] , \s_mux_signals[2][8][29] , 
        \s_mux_signals[2][8][28] , \s_mux_signals[2][8][27] , 
        \s_mux_signals[2][8][26] , \s_mux_signals[2][8][25] , 
        \s_mux_signals[2][8][24] , \s_mux_signals[2][8][23] , 
        \s_mux_signals[2][8][22] , \s_mux_signals[2][8][21] , 
        \s_mux_signals[2][8][20] , \s_mux_signals[2][8][19] , 
        \s_mux_signals[2][8][18] , \s_mux_signals[2][8][17] , 
        \s_mux_signals[2][8][16] , \s_mux_signals[2][8][15] , 
        \s_mux_signals[2][8][14] , \s_mux_signals[2][8][13] , 
        \s_mux_signals[2][8][12] , \s_mux_signals[2][8][11] , 
        \s_mux_signals[2][8][10] , \s_mux_signals[2][8][9] , 
        \s_mux_signals[2][8][8] , \s_mux_signals[2][8][7] , 
        \s_mux_signals[2][8][6] , \s_mux_signals[2][8][5] , 
        \s_mux_signals[2][8][4] , \s_mux_signals[2][8][3] , 
        \s_mux_signals[2][8][2] , \s_mux_signals[2][8][1] , 
        \s_mux_signals[2][8][0] }), .port1({\s_mux_signals[2][12][31] , 
        \s_mux_signals[2][12][30] , \s_mux_signals[2][12][29] , 
        \s_mux_signals[2][12][28] , \s_mux_signals[2][12][27] , 
        \s_mux_signals[2][12][26] , \s_mux_signals[2][12][25] , 
        \s_mux_signals[2][12][24] , \s_mux_signals[2][12][23] , 
        \s_mux_signals[2][12][22] , \s_mux_signals[2][12][21] , 
        \s_mux_signals[2][12][20] , \s_mux_signals[2][12][19] , 
        \s_mux_signals[2][12][18] , \s_mux_signals[2][12][17] , 
        \s_mux_signals[2][12][16] , \s_mux_signals[2][12][15] , 
        \s_mux_signals[2][12][14] , \s_mux_signals[2][12][13] , 
        \s_mux_signals[2][12][12] , \s_mux_signals[2][12][11] , 
        \s_mux_signals[2][12][10] , \s_mux_signals[2][12][9] , 
        \s_mux_signals[2][12][8] , \s_mux_signals[2][12][7] , 
        \s_mux_signals[2][12][6] , \s_mux_signals[2][12][5] , 
        \s_mux_signals[2][12][4] , \s_mux_signals[2][12][3] , 
        \s_mux_signals[2][12][2] , \s_mux_signals[2][12][1] , 
        \s_mux_signals[2][12][0] }), .sel(n26), .portY({
        \s_mux_signals[3][8][31] , \s_mux_signals[3][8][30] , 
        \s_mux_signals[3][8][29] , \s_mux_signals[3][8][28] , 
        \s_mux_signals[3][8][27] , \s_mux_signals[3][8][26] , 
        \s_mux_signals[3][8][25] , \s_mux_signals[3][8][24] , 
        \s_mux_signals[3][8][23] , \s_mux_signals[3][8][22] , 
        \s_mux_signals[3][8][21] , \s_mux_signals[3][8][20] , 
        \s_mux_signals[3][8][19] , \s_mux_signals[3][8][18] , 
        \s_mux_signals[3][8][17] , \s_mux_signals[3][8][16] , 
        \s_mux_signals[3][8][15] , \s_mux_signals[3][8][14] , 
        \s_mux_signals[3][8][13] , \s_mux_signals[3][8][12] , 
        \s_mux_signals[3][8][11] , \s_mux_signals[3][8][10] , 
        \s_mux_signals[3][8][9] , \s_mux_signals[3][8][8] , 
        \s_mux_signals[3][8][7] , \s_mux_signals[3][8][6] , 
        \s_mux_signals[3][8][5] , \s_mux_signals[3][8][4] , 
        \s_mux_signals[3][8][3] , \s_mux_signals[3][8][2] , 
        \s_mux_signals[3][8][1] , \s_mux_signals[3][8][0] }) );
  Mux_NBit_2x1_NBIT_IN32_95 MUX1_2_16 ( .port0({\s_mux_signals[2][16][31] , 
        \s_mux_signals[2][16][30] , \s_mux_signals[2][16][29] , 
        \s_mux_signals[2][16][28] , \s_mux_signals[2][16][27] , 
        \s_mux_signals[2][16][26] , \s_mux_signals[2][16][25] , 
        \s_mux_signals[2][16][24] , \s_mux_signals[2][16][23] , 
        \s_mux_signals[2][16][22] , \s_mux_signals[2][16][21] , 
        \s_mux_signals[2][16][20] , \s_mux_signals[2][16][19] , 
        \s_mux_signals[2][16][18] , \s_mux_signals[2][16][17] , 
        \s_mux_signals[2][16][16] , \s_mux_signals[2][16][15] , 
        \s_mux_signals[2][16][14] , \s_mux_signals[2][16][13] , 
        \s_mux_signals[2][16][12] , \s_mux_signals[2][16][11] , 
        \s_mux_signals[2][16][10] , \s_mux_signals[2][16][9] , 
        \s_mux_signals[2][16][8] , \s_mux_signals[2][16][7] , 
        \s_mux_signals[2][16][6] , \s_mux_signals[2][16][5] , 
        \s_mux_signals[2][16][4] , \s_mux_signals[2][16][3] , 
        \s_mux_signals[2][16][2] , \s_mux_signals[2][16][1] , 
        \s_mux_signals[2][16][0] }), .port1({\s_mux_signals[2][20][31] , 
        \s_mux_signals[2][20][30] , \s_mux_signals[2][20][29] , 
        \s_mux_signals[2][20][28] , \s_mux_signals[2][20][27] , 
        \s_mux_signals[2][20][26] , \s_mux_signals[2][20][25] , 
        \s_mux_signals[2][20][24] , \s_mux_signals[2][20][23] , 
        \s_mux_signals[2][20][22] , \s_mux_signals[2][20][21] , 
        \s_mux_signals[2][20][20] , \s_mux_signals[2][20][19] , 
        \s_mux_signals[2][20][18] , \s_mux_signals[2][20][17] , 
        \s_mux_signals[2][20][16] , \s_mux_signals[2][20][15] , 
        \s_mux_signals[2][20][14] , \s_mux_signals[2][20][13] , 
        \s_mux_signals[2][20][12] , \s_mux_signals[2][20][11] , 
        \s_mux_signals[2][20][10] , \s_mux_signals[2][20][9] , 
        \s_mux_signals[2][20][8] , \s_mux_signals[2][20][7] , 
        \s_mux_signals[2][20][6] , \s_mux_signals[2][20][5] , 
        \s_mux_signals[2][20][4] , \s_mux_signals[2][20][3] , 
        \s_mux_signals[2][20][2] , \s_mux_signals[2][20][1] , 
        \s_mux_signals[2][20][0] }), .sel(n26), .portY({
        \s_mux_signals[3][16][31] , \s_mux_signals[3][16][30] , 
        \s_mux_signals[3][16][29] , \s_mux_signals[3][16][28] , 
        \s_mux_signals[3][16][27] , \s_mux_signals[3][16][26] , 
        \s_mux_signals[3][16][25] , \s_mux_signals[3][16][24] , 
        \s_mux_signals[3][16][23] , \s_mux_signals[3][16][22] , 
        \s_mux_signals[3][16][21] , \s_mux_signals[3][16][20] , 
        \s_mux_signals[3][16][19] , \s_mux_signals[3][16][18] , 
        \s_mux_signals[3][16][17] , \s_mux_signals[3][16][16] , 
        \s_mux_signals[3][16][15] , \s_mux_signals[3][16][14] , 
        \s_mux_signals[3][16][13] , \s_mux_signals[3][16][12] , 
        \s_mux_signals[3][16][11] , \s_mux_signals[3][16][10] , 
        \s_mux_signals[3][16][9] , \s_mux_signals[3][16][8] , 
        \s_mux_signals[3][16][7] , \s_mux_signals[3][16][6] , 
        \s_mux_signals[3][16][5] , \s_mux_signals[3][16][4] , 
        \s_mux_signals[3][16][3] , \s_mux_signals[3][16][2] , 
        \s_mux_signals[3][16][1] , \s_mux_signals[3][16][0] }) );
  Mux_NBit_2x1_NBIT_IN32_94 MUX1_2_24 ( .port0({\s_mux_signals[2][24][31] , 
        \s_mux_signals[2][24][30] , \s_mux_signals[2][24][29] , 
        \s_mux_signals[2][24][28] , \s_mux_signals[2][24][27] , 
        \s_mux_signals[2][24][26] , \s_mux_signals[2][24][25] , 
        \s_mux_signals[2][24][24] , \s_mux_signals[2][24][23] , 
        \s_mux_signals[2][24][22] , \s_mux_signals[2][24][21] , 
        \s_mux_signals[2][24][20] , \s_mux_signals[2][24][19] , 
        \s_mux_signals[2][24][18] , \s_mux_signals[2][24][17] , 
        \s_mux_signals[2][24][16] , \s_mux_signals[2][24][15] , 
        \s_mux_signals[2][24][14] , \s_mux_signals[2][24][13] , 
        \s_mux_signals[2][24][12] , \s_mux_signals[2][24][11] , 
        \s_mux_signals[2][24][10] , \s_mux_signals[2][24][9] , 
        \s_mux_signals[2][24][8] , \s_mux_signals[2][24][7] , 
        \s_mux_signals[2][24][6] , \s_mux_signals[2][24][5] , 
        \s_mux_signals[2][24][4] , \s_mux_signals[2][24][3] , 
        \s_mux_signals[2][24][2] , \s_mux_signals[2][24][1] , 
        \s_mux_signals[2][24][0] }), .port1({\s_mux_signals[2][28][31] , 
        \s_mux_signals[2][28][30] , \s_mux_signals[2][28][29] , 
        \s_mux_signals[2][28][28] , \s_mux_signals[2][28][27] , 
        \s_mux_signals[2][28][26] , \s_mux_signals[2][28][25] , 
        \s_mux_signals[2][28][24] , \s_mux_signals[2][28][23] , 
        \s_mux_signals[2][28][22] , \s_mux_signals[2][28][21] , 
        \s_mux_signals[2][28][20] , \s_mux_signals[2][28][19] , 
        \s_mux_signals[2][28][18] , \s_mux_signals[2][28][17] , 
        \s_mux_signals[2][28][16] , \s_mux_signals[2][28][15] , 
        \s_mux_signals[2][28][14] , \s_mux_signals[2][28][13] , 
        \s_mux_signals[2][28][12] , \s_mux_signals[2][28][11] , 
        \s_mux_signals[2][28][10] , \s_mux_signals[2][28][9] , 
        \s_mux_signals[2][28][8] , \s_mux_signals[2][28][7] , 
        \s_mux_signals[2][28][6] , \s_mux_signals[2][28][5] , 
        \s_mux_signals[2][28][4] , \s_mux_signals[2][28][3] , 
        \s_mux_signals[2][28][2] , \s_mux_signals[2][28][1] , 
        \s_mux_signals[2][28][0] }), .sel(n26), .portY({
        \s_mux_signals[3][24][31] , \s_mux_signals[3][24][30] , 
        \s_mux_signals[3][24][29] , \s_mux_signals[3][24][28] , 
        \s_mux_signals[3][24][27] , \s_mux_signals[3][24][26] , 
        \s_mux_signals[3][24][25] , \s_mux_signals[3][24][24] , 
        \s_mux_signals[3][24][23] , \s_mux_signals[3][24][22] , 
        \s_mux_signals[3][24][21] , \s_mux_signals[3][24][20] , 
        \s_mux_signals[3][24][19] , \s_mux_signals[3][24][18] , 
        \s_mux_signals[3][24][17] , \s_mux_signals[3][24][16] , 
        \s_mux_signals[3][24][15] , \s_mux_signals[3][24][14] , 
        \s_mux_signals[3][24][13] , \s_mux_signals[3][24][12] , 
        \s_mux_signals[3][24][11] , \s_mux_signals[3][24][10] , 
        \s_mux_signals[3][24][9] , \s_mux_signals[3][24][8] , 
        \s_mux_signals[3][24][7] , \s_mux_signals[3][24][6] , 
        \s_mux_signals[3][24][5] , \s_mux_signals[3][24][4] , 
        \s_mux_signals[3][24][3] , \s_mux_signals[3][24][2] , 
        \s_mux_signals[3][24][1] , \s_mux_signals[3][24][0] }) );
  Mux_NBit_2x1_NBIT_IN32_93 MUX1_3_0 ( .port0({\s_mux_signals[3][0][31] , 
        \s_mux_signals[3][0][30] , \s_mux_signals[3][0][29] , 
        \s_mux_signals[3][0][28] , \s_mux_signals[3][0][27] , 
        \s_mux_signals[3][0][26] , \s_mux_signals[3][0][25] , 
        \s_mux_signals[3][0][24] , \s_mux_signals[3][0][23] , 
        \s_mux_signals[3][0][22] , \s_mux_signals[3][0][21] , 
        \s_mux_signals[3][0][20] , \s_mux_signals[3][0][19] , 
        \s_mux_signals[3][0][18] , \s_mux_signals[3][0][17] , 
        \s_mux_signals[3][0][16] , \s_mux_signals[3][0][15] , 
        \s_mux_signals[3][0][14] , \s_mux_signals[3][0][13] , 
        \s_mux_signals[3][0][12] , \s_mux_signals[3][0][11] , 
        \s_mux_signals[3][0][10] , \s_mux_signals[3][0][9] , 
        \s_mux_signals[3][0][8] , \s_mux_signals[3][0][7] , 
        \s_mux_signals[3][0][6] , \s_mux_signals[3][0][5] , 
        \s_mux_signals[3][0][4] , \s_mux_signals[3][0][3] , 
        \s_mux_signals[3][0][2] , \s_mux_signals[3][0][1] , 
        \s_mux_signals[3][0][0] }), .port1({\s_mux_signals[3][8][31] , 
        \s_mux_signals[3][8][30] , \s_mux_signals[3][8][29] , 
        \s_mux_signals[3][8][28] , \s_mux_signals[3][8][27] , 
        \s_mux_signals[3][8][26] , \s_mux_signals[3][8][25] , 
        \s_mux_signals[3][8][24] , \s_mux_signals[3][8][23] , 
        \s_mux_signals[3][8][22] , \s_mux_signals[3][8][21] , 
        \s_mux_signals[3][8][20] , \s_mux_signals[3][8][19] , 
        \s_mux_signals[3][8][18] , \s_mux_signals[3][8][17] , 
        \s_mux_signals[3][8][16] , \s_mux_signals[3][8][15] , 
        \s_mux_signals[3][8][14] , \s_mux_signals[3][8][13] , 
        \s_mux_signals[3][8][12] , \s_mux_signals[3][8][11] , 
        \s_mux_signals[3][8][10] , \s_mux_signals[3][8][9] , 
        \s_mux_signals[3][8][8] , \s_mux_signals[3][8][7] , 
        \s_mux_signals[3][8][6] , \s_mux_signals[3][8][5] , 
        \s_mux_signals[3][8][4] , \s_mux_signals[3][8][3] , 
        \s_mux_signals[3][8][2] , \s_mux_signals[3][8][1] , 
        \s_mux_signals[3][8][0] }), .sel(s_selmuxes_Fencoder_Tmuxes[3]), 
        .portY({\s_mux_signals[4][0][31] , \s_mux_signals[4][0][30] , 
        \s_mux_signals[4][0][29] , \s_mux_signals[4][0][28] , 
        \s_mux_signals[4][0][27] , \s_mux_signals[4][0][26] , 
        \s_mux_signals[4][0][25] , \s_mux_signals[4][0][24] , 
        \s_mux_signals[4][0][23] , \s_mux_signals[4][0][22] , 
        \s_mux_signals[4][0][21] , \s_mux_signals[4][0][20] , 
        \s_mux_signals[4][0][19] , \s_mux_signals[4][0][18] , 
        \s_mux_signals[4][0][17] , \s_mux_signals[4][0][16] , 
        \s_mux_signals[4][0][15] , \s_mux_signals[4][0][14] , 
        \s_mux_signals[4][0][13] , \s_mux_signals[4][0][12] , 
        \s_mux_signals[4][0][11] , \s_mux_signals[4][0][10] , 
        \s_mux_signals[4][0][9] , \s_mux_signals[4][0][8] , 
        \s_mux_signals[4][0][7] , \s_mux_signals[4][0][6] , 
        \s_mux_signals[4][0][5] , \s_mux_signals[4][0][4] , 
        \s_mux_signals[4][0][3] , \s_mux_signals[4][0][2] , 
        \s_mux_signals[4][0][1] , \s_mux_signals[4][0][0] }) );
  Mux_NBit_2x1_NBIT_IN32_92 MUX1_3_16 ( .port0({\s_mux_signals[3][16][31] , 
        \s_mux_signals[3][16][30] , \s_mux_signals[3][16][29] , 
        \s_mux_signals[3][16][28] , \s_mux_signals[3][16][27] , 
        \s_mux_signals[3][16][26] , \s_mux_signals[3][16][25] , 
        \s_mux_signals[3][16][24] , \s_mux_signals[3][16][23] , 
        \s_mux_signals[3][16][22] , \s_mux_signals[3][16][21] , 
        \s_mux_signals[3][16][20] , \s_mux_signals[3][16][19] , 
        \s_mux_signals[3][16][18] , \s_mux_signals[3][16][17] , 
        \s_mux_signals[3][16][16] , \s_mux_signals[3][16][15] , 
        \s_mux_signals[3][16][14] , \s_mux_signals[3][16][13] , 
        \s_mux_signals[3][16][12] , \s_mux_signals[3][16][11] , 
        \s_mux_signals[3][16][10] , \s_mux_signals[3][16][9] , 
        \s_mux_signals[3][16][8] , \s_mux_signals[3][16][7] , 
        \s_mux_signals[3][16][6] , \s_mux_signals[3][16][5] , 
        \s_mux_signals[3][16][4] , \s_mux_signals[3][16][3] , 
        \s_mux_signals[3][16][2] , \s_mux_signals[3][16][1] , 
        \s_mux_signals[3][16][0] }), .port1({\s_mux_signals[3][24][31] , 
        \s_mux_signals[3][24][30] , \s_mux_signals[3][24][29] , 
        \s_mux_signals[3][24][28] , \s_mux_signals[3][24][27] , 
        \s_mux_signals[3][24][26] , \s_mux_signals[3][24][25] , 
        \s_mux_signals[3][24][24] , \s_mux_signals[3][24][23] , 
        \s_mux_signals[3][24][22] , \s_mux_signals[3][24][21] , 
        \s_mux_signals[3][24][20] , \s_mux_signals[3][24][19] , 
        \s_mux_signals[3][24][18] , \s_mux_signals[3][24][17] , 
        \s_mux_signals[3][24][16] , \s_mux_signals[3][24][15] , 
        \s_mux_signals[3][24][14] , \s_mux_signals[3][24][13] , 
        \s_mux_signals[3][24][12] , \s_mux_signals[3][24][11] , 
        \s_mux_signals[3][24][10] , \s_mux_signals[3][24][9] , 
        \s_mux_signals[3][24][8] , \s_mux_signals[3][24][7] , 
        \s_mux_signals[3][24][6] , \s_mux_signals[3][24][5] , 
        \s_mux_signals[3][24][4] , \s_mux_signals[3][24][3] , 
        \s_mux_signals[3][24][2] , \s_mux_signals[3][24][1] , 
        \s_mux_signals[3][24][0] }), .sel(s_selmuxes_Fencoder_Tmuxes[3]), 
        .portY({\s_mux_signals[4][16][31] , \s_mux_signals[4][16][30] , 
        \s_mux_signals[4][16][29] , \s_mux_signals[4][16][28] , 
        \s_mux_signals[4][16][27] , \s_mux_signals[4][16][26] , 
        \s_mux_signals[4][16][25] , \s_mux_signals[4][16][24] , 
        \s_mux_signals[4][16][23] , \s_mux_signals[4][16][22] , 
        \s_mux_signals[4][16][21] , \s_mux_signals[4][16][20] , 
        \s_mux_signals[4][16][19] , \s_mux_signals[4][16][18] , 
        \s_mux_signals[4][16][17] , \s_mux_signals[4][16][16] , 
        \s_mux_signals[4][16][15] , \s_mux_signals[4][16][14] , 
        \s_mux_signals[4][16][13] , \s_mux_signals[4][16][12] , 
        \s_mux_signals[4][16][11] , \s_mux_signals[4][16][10] , 
        \s_mux_signals[4][16][9] , \s_mux_signals[4][16][8] , 
        \s_mux_signals[4][16][7] , \s_mux_signals[4][16][6] , 
        \s_mux_signals[4][16][5] , \s_mux_signals[4][16][4] , 
        \s_mux_signals[4][16][3] , \s_mux_signals[4][16][2] , 
        \s_mux_signals[4][16][1] , \s_mux_signals[4][16][0] }) );
  Mux_NBit_2x1_NBIT_IN32_91 MUX1_4_0 ( .port0({\s_mux_signals[4][0][31] , 
        \s_mux_signals[4][0][30] , \s_mux_signals[4][0][29] , 
        \s_mux_signals[4][0][28] , \s_mux_signals[4][0][27] , 
        \s_mux_signals[4][0][26] , \s_mux_signals[4][0][25] , 
        \s_mux_signals[4][0][24] , \s_mux_signals[4][0][23] , 
        \s_mux_signals[4][0][22] , \s_mux_signals[4][0][21] , 
        \s_mux_signals[4][0][20] , \s_mux_signals[4][0][19] , 
        \s_mux_signals[4][0][18] , \s_mux_signals[4][0][17] , 
        \s_mux_signals[4][0][16] , \s_mux_signals[4][0][15] , 
        \s_mux_signals[4][0][14] , \s_mux_signals[4][0][13] , 
        \s_mux_signals[4][0][12] , \s_mux_signals[4][0][11] , 
        \s_mux_signals[4][0][10] , \s_mux_signals[4][0][9] , 
        \s_mux_signals[4][0][8] , \s_mux_signals[4][0][7] , 
        \s_mux_signals[4][0][6] , \s_mux_signals[4][0][5] , 
        \s_mux_signals[4][0][4] , \s_mux_signals[4][0][3] , 
        \s_mux_signals[4][0][2] , \s_mux_signals[4][0][1] , 
        \s_mux_signals[4][0][0] }), .port1({\s_mux_signals[4][16][31] , 
        \s_mux_signals[4][16][30] , \s_mux_signals[4][16][29] , 
        \s_mux_signals[4][16][28] , \s_mux_signals[4][16][27] , 
        \s_mux_signals[4][16][26] , \s_mux_signals[4][16][25] , 
        \s_mux_signals[4][16][24] , \s_mux_signals[4][16][23] , 
        \s_mux_signals[4][16][22] , \s_mux_signals[4][16][21] , 
        \s_mux_signals[4][16][20] , \s_mux_signals[4][16][19] , 
        \s_mux_signals[4][16][18] , \s_mux_signals[4][16][17] , 
        \s_mux_signals[4][16][16] , \s_mux_signals[4][16][15] , 
        \s_mux_signals[4][16][14] , \s_mux_signals[4][16][13] , 
        \s_mux_signals[4][16][12] , \s_mux_signals[4][16][11] , 
        \s_mux_signals[4][16][10] , \s_mux_signals[4][16][9] , 
        \s_mux_signals[4][16][8] , \s_mux_signals[4][16][7] , 
        \s_mux_signals[4][16][6] , \s_mux_signals[4][16][5] , 
        \s_mux_signals[4][16][4] , \s_mux_signals[4][16][3] , 
        \s_mux_signals[4][16][2] , \s_mux_signals[4][16][1] , 
        \s_mux_signals[4][16][0] }), .sel(s_selmuxes_Fencoder_Tmuxes[4]), 
        .portY({\s_mux_signals[5][0][31] , \s_mux_signals[5][0][30] , 
        \s_mux_signals[5][0][29] , \s_mux_signals[5][0][28] , 
        \s_mux_signals[5][0][27] , \s_mux_signals[5][0][26] , 
        \s_mux_signals[5][0][25] , \s_mux_signals[5][0][24] , 
        \s_mux_signals[5][0][23] , \s_mux_signals[5][0][22] , 
        \s_mux_signals[5][0][21] , \s_mux_signals[5][0][20] , 
        \s_mux_signals[5][0][19] , \s_mux_signals[5][0][18] , 
        \s_mux_signals[5][0][17] , \s_mux_signals[5][0][16] , 
        \s_mux_signals[5][0][15] , \s_mux_signals[5][0][14] , 
        \s_mux_signals[5][0][13] , \s_mux_signals[5][0][12] , 
        \s_mux_signals[5][0][11] , \s_mux_signals[5][0][10] , 
        \s_mux_signals[5][0][9] , \s_mux_signals[5][0][8] , 
        \s_mux_signals[5][0][7] , \s_mux_signals[5][0][6] , 
        \s_mux_signals[5][0][5] , \s_mux_signals[5][0][4] , 
        \s_mux_signals[5][0][3] , \s_mux_signals[5][0][2] , 
        \s_mux_signals[5][0][1] , \s_mux_signals[5][0][0] }) );
  Mux_NBit_2x1_NBIT_IN32_90 MuxTargOut ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0}), .port1({\s_mux_signals[5][0][31] , 
        \s_mux_signals[5][0][30] , \s_mux_signals[5][0][29] , 
        \s_mux_signals[5][0][28] , \s_mux_signals[5][0][27] , 
        \s_mux_signals[5][0][26] , \s_mux_signals[5][0][25] , 
        \s_mux_signals[5][0][24] , \s_mux_signals[5][0][23] , 
        \s_mux_signals[5][0][22] , \s_mux_signals[5][0][21] , 
        \s_mux_signals[5][0][20] , \s_mux_signals[5][0][19] , 
        \s_mux_signals[5][0][18] , \s_mux_signals[5][0][17] , 
        \s_mux_signals[5][0][16] , \s_mux_signals[5][0][15] , 
        \s_mux_signals[5][0][14] , \s_mux_signals[5][0][13] , 
        \s_mux_signals[5][0][12] , \s_mux_signals[5][0][11] , 
        \s_mux_signals[5][0][10] , \s_mux_signals[5][0][9] , 
        \s_mux_signals[5][0][8] , \s_mux_signals[5][0][7] , 
        \s_mux_signals[5][0][6] , \s_mux_signals[5][0][5] , 
        \s_mux_signals[5][0][4] , \s_mux_signals[5][0][3] , 
        \s_mux_signals[5][0][2] , \s_mux_signals[5][0][1] , 
        \s_mux_signals[5][0][0] }), .sel(s_HIT_miss), .portY(
        BTB_target_prediction) );
  BUF_X2 U3 ( .A(BTB_target_From_DE[31]), .Z(n125) );
  BUF_X1 U4 ( .A(BTB_target_From_DE[19]), .Z(n87) );
  BUF_X1 U5 ( .A(BTB_target_From_DE[19]), .Z(n88) );
  BUF_X1 U6 ( .A(BTB_target_From_DE[20]), .Z(n90) );
  BUF_X1 U7 ( .A(BTB_target_From_DE[21]), .Z(n93) );
  BUF_X1 U8 ( .A(BTB_target_From_DE[22]), .Z(n96) );
  BUF_X1 U9 ( .A(BTB_target_From_DE[23]), .Z(n99) );
  BUF_X1 U10 ( .A(BTB_target_From_DE[24]), .Z(n102) );
  BUF_X1 U11 ( .A(BTB_target_From_DE[20]), .Z(n91) );
  BUF_X1 U12 ( .A(BTB_target_From_DE[21]), .Z(n94) );
  BUF_X1 U13 ( .A(BTB_target_From_DE[22]), .Z(n97) );
  BUF_X1 U14 ( .A(BTB_target_From_DE[23]), .Z(n100) );
  BUF_X1 U15 ( .A(BTB_target_From_DE[24]), .Z(n103) );
  BUF_X1 U16 ( .A(BTB_target_From_DE[25]), .Z(n107) );
  BUF_X1 U17 ( .A(BTB_target_From_DE[26]), .Z(n110) );
  BUF_X1 U18 ( .A(BTB_target_From_DE[27]), .Z(n113) );
  BUF_X1 U19 ( .A(BTB_target_From_DE[28]), .Z(n116) );
  BUF_X1 U20 ( .A(BTB_target_From_DE[29]), .Z(n119) );
  BUF_X1 U21 ( .A(BTB_target_From_DE[30]), .Z(n122) );
  BUF_X1 U22 ( .A(n326), .Z(n333) );
  BUF_X1 U23 ( .A(n326), .Z(n332) );
  BUF_X1 U24 ( .A(n326), .Z(n331) );
  BUF_X1 U25 ( .A(n325), .Z(n330) );
  BUF_X1 U26 ( .A(n325), .Z(n329) );
  BUF_X1 U27 ( .A(n325), .Z(n328) );
  BUF_X1 U28 ( .A(n15), .Z(n17) );
  BUF_X1 U29 ( .A(n15), .Z(n18) );
  BUF_X1 U30 ( .A(n15), .Z(n19) );
  BUF_X1 U31 ( .A(n16), .Z(n20) );
  BUF_X1 U32 ( .A(n16), .Z(n21) );
  BUF_X1 U33 ( .A(n16), .Z(n22) );
  INV_X1 U34 ( .A(n8), .ZN(n324) );
  BUF_X1 U35 ( .A(n1), .Z(n15) );
  BUF_X1 U36 ( .A(n1), .Z(n16) );
  BUF_X2 U37 ( .A(BTB_target_From_DE[31]), .Z(n123) );
  BUF_X2 U38 ( .A(BTB_target_From_DE[31]), .Z(n124) );
  BUF_X2 U39 ( .A(BTB_target_From_DE[30]), .Z(n120) );
  BUF_X2 U40 ( .A(BTB_target_From_DE[30]), .Z(n121) );
  BUF_X2 U41 ( .A(BTB_target_From_DE[29]), .Z(n117) );
  BUF_X2 U42 ( .A(BTB_target_From_DE[29]), .Z(n118) );
  BUF_X2 U43 ( .A(BTB_target_From_DE[28]), .Z(n114) );
  BUF_X2 U44 ( .A(BTB_target_From_DE[28]), .Z(n115) );
  BUF_X2 U45 ( .A(BTB_target_From_DE[27]), .Z(n111) );
  BUF_X2 U46 ( .A(BTB_target_From_DE[27]), .Z(n112) );
  BUF_X2 U47 ( .A(BTB_target_From_DE[26]), .Z(n108) );
  BUF_X2 U48 ( .A(BTB_target_From_DE[26]), .Z(n109) );
  BUF_X1 U49 ( .A(BTB_branch_taken), .Z(n27) );
  BUF_X1 U50 ( .A(BTB_branch_taken), .Z(n28) );
  BUF_X1 U51 ( .A(BTB_branch_taken), .Z(n29) );
  BUF_X2 U52 ( .A(BTB_target_From_DE[25]), .Z(n105) );
  BUF_X2 U53 ( .A(BTB_target_From_DE[25]), .Z(n106) );
  BUF_X1 U54 ( .A(BTB_target_From_DE[18]), .Z(n84) );
  BUF_X1 U55 ( .A(BTB_target_From_DE[18]), .Z(n85) );
  BUF_X1 U56 ( .A(BTB_target_From_DE[13]), .Z(n69) );
  BUF_X1 U57 ( .A(BTB_target_From_DE[14]), .Z(n72) );
  BUF_X1 U58 ( .A(BTB_target_From_DE[13]), .Z(n70) );
  BUF_X1 U59 ( .A(BTB_target_From_DE[14]), .Z(n73) );
  BUF_X1 U60 ( .A(BTB_target_From_DE[17]), .Z(n81) );
  BUF_X1 U61 ( .A(BTB_target_From_DE[17]), .Z(n82) );
  BUF_X1 U62 ( .A(BTB_target_From_DE[16]), .Z(n78) );
  BUF_X1 U63 ( .A(BTB_target_From_DE[16]), .Z(n79) );
  BUF_X1 U64 ( .A(BTB_target_From_DE[15]), .Z(n75) );
  BUF_X1 U65 ( .A(BTB_target_From_DE[15]), .Z(n76) );
  BUF_X1 U66 ( .A(BTB_target_From_DE[4]), .Z(n42) );
  BUF_X1 U67 ( .A(BTB_target_From_DE[5]), .Z(n45) );
  BUF_X1 U68 ( .A(BTB_target_From_DE[6]), .Z(n48) );
  BUF_X1 U69 ( .A(BTB_target_From_DE[7]), .Z(n51) );
  BUF_X1 U70 ( .A(BTB_target_From_DE[8]), .Z(n54) );
  BUF_X1 U71 ( .A(BTB_target_From_DE[9]), .Z(n57) );
  BUF_X1 U72 ( .A(BTB_target_From_DE[10]), .Z(n60) );
  BUF_X1 U73 ( .A(BTB_target_From_DE[11]), .Z(n63) );
  BUF_X1 U74 ( .A(BTB_target_From_DE[12]), .Z(n66) );
  BUF_X1 U75 ( .A(BTB_target_From_DE[4]), .Z(n43) );
  BUF_X1 U76 ( .A(BTB_target_From_DE[5]), .Z(n46) );
  BUF_X1 U77 ( .A(BTB_target_From_DE[6]), .Z(n49) );
  BUF_X1 U78 ( .A(BTB_target_From_DE[7]), .Z(n52) );
  BUF_X1 U79 ( .A(BTB_target_From_DE[8]), .Z(n55) );
  BUF_X1 U80 ( .A(BTB_target_From_DE[9]), .Z(n58) );
  BUF_X1 U81 ( .A(BTB_target_From_DE[10]), .Z(n61) );
  BUF_X1 U82 ( .A(BTB_target_From_DE[11]), .Z(n64) );
  BUF_X1 U83 ( .A(BTB_target_From_DE[12]), .Z(n67) );
  BUF_X1 U84 ( .A(BTB_target_From_DE[24]), .Z(n104) );
  BUF_X1 U85 ( .A(BTB_target_From_DE[23]), .Z(n101) );
  BUF_X1 U86 ( .A(BTB_target_From_DE[22]), .Z(n98) );
  BUF_X1 U87 ( .A(BTB_target_From_DE[21]), .Z(n95) );
  BUF_X1 U88 ( .A(BTB_target_From_DE[20]), .Z(n92) );
  BUF_X1 U89 ( .A(BTB_target_From_DE[19]), .Z(n89) );
  BUF_X1 U90 ( .A(BTB_target_From_DE[18]), .Z(n86) );
  BUF_X1 U91 ( .A(BTB_target_From_DE[13]), .Z(n71) );
  BUF_X1 U92 ( .A(BTB_target_From_DE[14]), .Z(n74) );
  BUF_X1 U93 ( .A(BTB_target_From_DE[17]), .Z(n83) );
  BUF_X1 U94 ( .A(BTB_target_From_DE[16]), .Z(n80) );
  BUF_X1 U95 ( .A(BTB_target_From_DE[15]), .Z(n77) );
  BUF_X1 U96 ( .A(BTB_target_From_DE[4]), .Z(n44) );
  BUF_X1 U97 ( .A(BTB_target_From_DE[5]), .Z(n47) );
  BUF_X1 U98 ( .A(BTB_target_From_DE[6]), .Z(n50) );
  BUF_X1 U99 ( .A(BTB_target_From_DE[7]), .Z(n53) );
  BUF_X1 U100 ( .A(BTB_target_From_DE[8]), .Z(n56) );
  BUF_X1 U101 ( .A(BTB_target_From_DE[9]), .Z(n59) );
  BUF_X1 U102 ( .A(BTB_target_From_DE[10]), .Z(n62) );
  BUF_X1 U103 ( .A(BTB_target_From_DE[11]), .Z(n65) );
  BUF_X1 U104 ( .A(BTB_target_From_DE[12]), .Z(n68) );
  BUF_X1 U105 ( .A(BTB_PC_From_IF[20]), .Z(n282) );
  BUF_X1 U106 ( .A(BTB_PC_From_IF[21]), .Z(n285) );
  BUF_X1 U107 ( .A(BTB_PC_From_IF[22]), .Z(n288) );
  BUF_X1 U108 ( .A(BTB_PC_From_IF[23]), .Z(n291) );
  BUF_X1 U109 ( .A(BTB_PC_From_IF[17]), .Z(n273) );
  BUF_X1 U110 ( .A(BTB_PC_From_IF[18]), .Z(n276) );
  BUF_X1 U111 ( .A(BTB_PC_From_IF[19]), .Z(n279) );
  BUF_X1 U112 ( .A(BTB_PC_From_IF[1]), .Z(n225) );
  BUF_X1 U113 ( .A(BTB_PC_From_IF[13]), .Z(n261) );
  BUF_X1 U114 ( .A(BTB_PC_From_IF[14]), .Z(n264) );
  BUF_X1 U115 ( .A(BTB_PC_From_IF[15]), .Z(n267) );
  BUF_X1 U116 ( .A(BTB_PC_From_IF[16]), .Z(n270) );
  BUF_X1 U117 ( .A(BTB_PC_From_IF[0]), .Z(n222) );
  BUF_X1 U118 ( .A(BTB_PC_From_IF[10]), .Z(n252) );
  BUF_X1 U119 ( .A(BTB_PC_From_IF[11]), .Z(n255) );
  BUF_X1 U120 ( .A(BTB_PC_From_IF[12]), .Z(n258) );
  BUF_X1 U121 ( .A(BTB_PC_From_IF[6]), .Z(n240) );
  BUF_X1 U122 ( .A(BTB_PC_From_IF[7]), .Z(n243) );
  BUF_X1 U123 ( .A(BTB_PC_From_IF[8]), .Z(n246) );
  BUF_X1 U124 ( .A(BTB_PC_From_IF[9]), .Z(n249) );
  BUF_X1 U125 ( .A(BTB_PC_From_IF[3]), .Z(n231) );
  BUF_X1 U126 ( .A(BTB_PC_From_IF[31]), .Z(n315) );
  BUF_X1 U127 ( .A(BTB_PC_From_IF[4]), .Z(n234) );
  BUF_X1 U128 ( .A(BTB_PC_From_IF[5]), .Z(n237) );
  BUF_X1 U129 ( .A(BTB_PC_From_IF[2]), .Z(n228) );
  BUF_X1 U130 ( .A(BTB_PC_From_IF[28]), .Z(n306) );
  BUF_X1 U131 ( .A(BTB_PC_From_IF[29]), .Z(n309) );
  BUF_X1 U132 ( .A(BTB_PC_From_IF[30]), .Z(n312) );
  BUF_X1 U133 ( .A(BTB_PC_From_IF[24]), .Z(n294) );
  BUF_X1 U134 ( .A(BTB_PC_From_IF[25]), .Z(n297) );
  BUF_X1 U135 ( .A(BTB_PC_From_IF[26]), .Z(n300) );
  BUF_X1 U136 ( .A(BTB_PC_From_IF[27]), .Z(n303) );
  BUF_X1 U137 ( .A(BTB_PC_From_IF[20]), .Z(n283) );
  BUF_X1 U138 ( .A(BTB_PC_From_IF[21]), .Z(n286) );
  BUF_X1 U139 ( .A(BTB_PC_From_IF[22]), .Z(n289) );
  BUF_X1 U140 ( .A(BTB_PC_From_IF[23]), .Z(n292) );
  BUF_X1 U141 ( .A(BTB_PC_From_IF[17]), .Z(n274) );
  BUF_X1 U142 ( .A(BTB_PC_From_IF[18]), .Z(n277) );
  BUF_X1 U143 ( .A(BTB_PC_From_IF[19]), .Z(n280) );
  BUF_X1 U144 ( .A(BTB_PC_From_IF[1]), .Z(n226) );
  BUF_X1 U145 ( .A(BTB_PC_From_IF[13]), .Z(n262) );
  BUF_X1 U146 ( .A(BTB_PC_From_IF[14]), .Z(n265) );
  BUF_X1 U147 ( .A(BTB_PC_From_IF[15]), .Z(n268) );
  BUF_X1 U148 ( .A(BTB_PC_From_IF[16]), .Z(n271) );
  BUF_X1 U149 ( .A(BTB_PC_From_IF[0]), .Z(n223) );
  BUF_X1 U150 ( .A(BTB_PC_From_IF[10]), .Z(n253) );
  BUF_X1 U151 ( .A(BTB_PC_From_IF[11]), .Z(n256) );
  BUF_X1 U152 ( .A(BTB_PC_From_IF[12]), .Z(n259) );
  BUF_X1 U153 ( .A(BTB_PC_From_IF[6]), .Z(n241) );
  BUF_X1 U154 ( .A(BTB_PC_From_IF[7]), .Z(n244) );
  BUF_X1 U155 ( .A(BTB_PC_From_IF[8]), .Z(n247) );
  BUF_X1 U156 ( .A(BTB_PC_From_IF[9]), .Z(n250) );
  BUF_X1 U157 ( .A(BTB_PC_From_IF[3]), .Z(n232) );
  BUF_X1 U158 ( .A(BTB_PC_From_IF[4]), .Z(n235) );
  BUF_X1 U159 ( .A(BTB_PC_From_IF[31]), .Z(n316) );
  BUF_X1 U160 ( .A(BTB_PC_From_IF[5]), .Z(n238) );
  BUF_X1 U161 ( .A(BTB_PC_From_IF[2]), .Z(n229) );
  BUF_X1 U162 ( .A(BTB_PC_From_IF[28]), .Z(n307) );
  BUF_X1 U163 ( .A(BTB_PC_From_IF[29]), .Z(n310) );
  BUF_X1 U164 ( .A(BTB_PC_From_IF[30]), .Z(n313) );
  BUF_X1 U165 ( .A(BTB_PC_From_IF[24]), .Z(n295) );
  BUF_X1 U166 ( .A(BTB_PC_From_IF[25]), .Z(n298) );
  BUF_X1 U167 ( .A(BTB_PC_From_IF[26]), .Z(n301) );
  BUF_X1 U168 ( .A(BTB_PC_From_IF[27]), .Z(n304) );
  BUF_X1 U169 ( .A(BTB_target_From_DE[1]), .Z(n33) );
  BUF_X1 U170 ( .A(BTB_target_From_DE[2]), .Z(n36) );
  BUF_X1 U171 ( .A(BTB_target_From_DE[3]), .Z(n39) );
  BUF_X1 U172 ( .A(BTB_target_From_DE[1]), .Z(n34) );
  BUF_X1 U173 ( .A(BTB_target_From_DE[2]), .Z(n37) );
  BUF_X1 U174 ( .A(BTB_target_From_DE[3]), .Z(n40) );
  BUF_X1 U175 ( .A(BTB_target_From_DE[1]), .Z(n35) );
  BUF_X1 U176 ( .A(BTB_target_From_DE[2]), .Z(n38) );
  BUF_X1 U177 ( .A(BTB_target_From_DE[3]), .Z(n41) );
  BUF_X1 U178 ( .A(BTB_PC_From_IF[20]), .Z(n284) );
  BUF_X1 U179 ( .A(BTB_PC_From_IF[21]), .Z(n287) );
  BUF_X1 U180 ( .A(BTB_PC_From_IF[22]), .Z(n290) );
  BUF_X1 U181 ( .A(BTB_PC_From_IF[23]), .Z(n293) );
  BUF_X1 U182 ( .A(BTB_PC_From_IF[17]), .Z(n275) );
  BUF_X1 U183 ( .A(BTB_PC_From_IF[18]), .Z(n278) );
  BUF_X1 U184 ( .A(BTB_PC_From_IF[19]), .Z(n281) );
  BUF_X1 U185 ( .A(BTB_PC_From_IF[1]), .Z(n227) );
  BUF_X1 U186 ( .A(BTB_PC_From_IF[13]), .Z(n263) );
  BUF_X1 U187 ( .A(BTB_PC_From_IF[14]), .Z(n266) );
  BUF_X1 U188 ( .A(BTB_PC_From_IF[15]), .Z(n269) );
  BUF_X1 U189 ( .A(BTB_PC_From_IF[16]), .Z(n272) );
  BUF_X1 U190 ( .A(BTB_PC_From_IF[0]), .Z(n224) );
  BUF_X1 U191 ( .A(BTB_PC_From_IF[10]), .Z(n254) );
  BUF_X1 U192 ( .A(BTB_PC_From_IF[11]), .Z(n257) );
  BUF_X1 U193 ( .A(BTB_PC_From_IF[12]), .Z(n260) );
  BUF_X1 U194 ( .A(BTB_PC_From_IF[6]), .Z(n242) );
  BUF_X1 U195 ( .A(BTB_PC_From_IF[7]), .Z(n245) );
  BUF_X1 U196 ( .A(BTB_PC_From_IF[8]), .Z(n248) );
  BUF_X1 U197 ( .A(BTB_PC_From_IF[9]), .Z(n251) );
  BUF_X1 U198 ( .A(BTB_PC_From_IF[3]), .Z(n233) );
  BUF_X1 U199 ( .A(BTB_PC_From_IF[31]), .Z(n317) );
  BUF_X1 U200 ( .A(BTB_PC_From_IF[4]), .Z(n236) );
  BUF_X1 U201 ( .A(BTB_PC_From_IF[5]), .Z(n239) );
  BUF_X1 U202 ( .A(BTB_PC_From_IF[2]), .Z(n230) );
  BUF_X1 U203 ( .A(BTB_PC_From_IF[28]), .Z(n308) );
  BUF_X1 U204 ( .A(BTB_PC_From_IF[29]), .Z(n311) );
  BUF_X1 U205 ( .A(BTB_PC_From_IF[30]), .Z(n314) );
  BUF_X1 U206 ( .A(BTB_PC_From_IF[24]), .Z(n296) );
  BUF_X1 U207 ( .A(BTB_PC_From_IF[25]), .Z(n299) );
  BUF_X1 U208 ( .A(BTB_PC_From_IF[26]), .Z(n302) );
  BUF_X1 U209 ( .A(BTB_PC_From_IF[27]), .Z(n305) );
  NOR2_X1 U210 ( .A1(BTB_restore), .A2(n324), .ZN(n1) );
  BUF_X2 U211 ( .A(n327), .Z(n334) );
  BUF_X1 U212 ( .A(n327), .Z(n335) );
  BUF_X1 U213 ( .A(BTB_PC_From_DE[2]), .Z(n132) );
  BUF_X1 U214 ( .A(BTB_PC_From_DE[3]), .Z(n135) );
  BUF_X1 U215 ( .A(BTB_PC_From_DE[4]), .Z(n138) );
  BUF_X1 U216 ( .A(BTB_PC_From_DE[5]), .Z(n141) );
  BUF_X1 U217 ( .A(BTB_PC_From_DE[6]), .Z(n144) );
  BUF_X1 U218 ( .A(BTB_PC_From_DE[7]), .Z(n147) );
  BUF_X1 U219 ( .A(BTB_PC_From_DE[30]), .Z(n216) );
  BUF_X1 U220 ( .A(BTB_PC_From_DE[31]), .Z(n219) );
  BUF_X1 U221 ( .A(BTB_PC_From_DE[2]), .Z(n133) );
  BUF_X1 U222 ( .A(BTB_PC_From_DE[3]), .Z(n136) );
  BUF_X1 U223 ( .A(BTB_PC_From_DE[4]), .Z(n139) );
  BUF_X1 U224 ( .A(BTB_PC_From_DE[5]), .Z(n142) );
  BUF_X1 U225 ( .A(BTB_PC_From_DE[6]), .Z(n145) );
  BUF_X1 U226 ( .A(BTB_PC_From_DE[7]), .Z(n148) );
  BUF_X1 U227 ( .A(BTB_PC_From_DE[30]), .Z(n217) );
  BUF_X1 U228 ( .A(BTB_PC_From_DE[31]), .Z(n220) );
  BUF_X1 U229 ( .A(BTB_PC_From_DE[0]), .Z(n126) );
  BUF_X1 U230 ( .A(BTB_PC_From_DE[1]), .Z(n129) );
  BUF_X1 U231 ( .A(BTB_PC_From_DE[8]), .Z(n150) );
  BUF_X1 U232 ( .A(BTB_PC_From_DE[9]), .Z(n153) );
  BUF_X1 U233 ( .A(BTB_PC_From_DE[10]), .Z(n156) );
  BUF_X1 U234 ( .A(BTB_PC_From_DE[11]), .Z(n159) );
  BUF_X1 U235 ( .A(BTB_PC_From_DE[12]), .Z(n162) );
  BUF_X1 U236 ( .A(BTB_PC_From_DE[13]), .Z(n165) );
  BUF_X1 U237 ( .A(BTB_PC_From_DE[14]), .Z(n168) );
  BUF_X1 U238 ( .A(BTB_PC_From_DE[15]), .Z(n171) );
  BUF_X1 U239 ( .A(BTB_PC_From_DE[16]), .Z(n174) );
  BUF_X1 U240 ( .A(BTB_PC_From_DE[17]), .Z(n177) );
  BUF_X1 U241 ( .A(BTB_PC_From_DE[18]), .Z(n180) );
  BUF_X1 U242 ( .A(BTB_PC_From_DE[19]), .Z(n183) );
  BUF_X1 U243 ( .A(BTB_PC_From_DE[20]), .Z(n186) );
  BUF_X1 U244 ( .A(BTB_PC_From_DE[21]), .Z(n189) );
  BUF_X1 U245 ( .A(BTB_PC_From_DE[22]), .Z(n192) );
  BUF_X1 U246 ( .A(BTB_PC_From_DE[23]), .Z(n195) );
  BUF_X1 U247 ( .A(BTB_PC_From_DE[24]), .Z(n198) );
  BUF_X1 U248 ( .A(BTB_PC_From_DE[25]), .Z(n201) );
  BUF_X1 U249 ( .A(BTB_PC_From_DE[26]), .Z(n204) );
  BUF_X1 U250 ( .A(BTB_PC_From_DE[27]), .Z(n207) );
  BUF_X1 U251 ( .A(BTB_PC_From_DE[28]), .Z(n210) );
  BUF_X1 U252 ( .A(BTB_PC_From_DE[29]), .Z(n213) );
  BUF_X1 U253 ( .A(BTB_PC_From_DE[0]), .Z(n127) );
  BUF_X1 U254 ( .A(BTB_PC_From_DE[1]), .Z(n130) );
  BUF_X1 U255 ( .A(BTB_PC_From_DE[8]), .Z(n151) );
  BUF_X1 U256 ( .A(BTB_PC_From_DE[9]), .Z(n154) );
  BUF_X1 U257 ( .A(BTB_PC_From_DE[10]), .Z(n157) );
  BUF_X1 U258 ( .A(BTB_PC_From_DE[11]), .Z(n160) );
  BUF_X1 U259 ( .A(BTB_PC_From_DE[12]), .Z(n163) );
  BUF_X1 U260 ( .A(BTB_PC_From_DE[13]), .Z(n166) );
  BUF_X1 U261 ( .A(BTB_PC_From_DE[14]), .Z(n169) );
  BUF_X1 U262 ( .A(BTB_PC_From_DE[15]), .Z(n172) );
  BUF_X1 U263 ( .A(BTB_PC_From_DE[16]), .Z(n175) );
  BUF_X1 U264 ( .A(BTB_PC_From_DE[17]), .Z(n178) );
  BUF_X1 U265 ( .A(BTB_PC_From_DE[18]), .Z(n181) );
  BUF_X1 U266 ( .A(BTB_PC_From_DE[19]), .Z(n184) );
  BUF_X1 U267 ( .A(BTB_PC_From_DE[20]), .Z(n187) );
  BUF_X1 U268 ( .A(BTB_PC_From_DE[21]), .Z(n190) );
  BUF_X1 U269 ( .A(BTB_PC_From_DE[22]), .Z(n193) );
  BUF_X1 U270 ( .A(BTB_PC_From_DE[23]), .Z(n196) );
  BUF_X1 U271 ( .A(BTB_PC_From_DE[24]), .Z(n199) );
  BUF_X1 U272 ( .A(BTB_PC_From_DE[25]), .Z(n202) );
  BUF_X1 U273 ( .A(BTB_PC_From_DE[26]), .Z(n205) );
  BUF_X1 U274 ( .A(BTB_PC_From_DE[27]), .Z(n208) );
  BUF_X1 U275 ( .A(BTB_PC_From_DE[28]), .Z(n211) );
  BUF_X1 U276 ( .A(BTB_PC_From_DE[29]), .Z(n214) );
  BUF_X1 U277 ( .A(BTB_target_From_DE[0]), .Z(n30) );
  BUF_X1 U278 ( .A(BTB_target_From_DE[0]), .Z(n31) );
  BUF_X1 U279 ( .A(BTB_PC_From_DE[2]), .Z(n134) );
  BUF_X1 U280 ( .A(BTB_PC_From_DE[3]), .Z(n137) );
  BUF_X1 U281 ( .A(BTB_PC_From_DE[4]), .Z(n140) );
  BUF_X1 U282 ( .A(BTB_PC_From_DE[5]), .Z(n143) );
  BUF_X1 U283 ( .A(BTB_PC_From_DE[6]), .Z(n146) );
  BUF_X1 U284 ( .A(BTB_PC_From_DE[7]), .Z(n149) );
  BUF_X1 U285 ( .A(BTB_PC_From_DE[30]), .Z(n218) );
  BUF_X1 U286 ( .A(BTB_PC_From_DE[31]), .Z(n221) );
  BUF_X1 U287 ( .A(BTB_PC_From_DE[0]), .Z(n128) );
  BUF_X1 U288 ( .A(BTB_PC_From_DE[1]), .Z(n131) );
  BUF_X1 U289 ( .A(BTB_PC_From_DE[8]), .Z(n152) );
  BUF_X1 U290 ( .A(BTB_PC_From_DE[9]), .Z(n155) );
  BUF_X1 U291 ( .A(BTB_PC_From_DE[10]), .Z(n158) );
  BUF_X1 U292 ( .A(BTB_PC_From_DE[11]), .Z(n161) );
  BUF_X1 U293 ( .A(BTB_PC_From_DE[12]), .Z(n164) );
  BUF_X1 U294 ( .A(BTB_PC_From_DE[13]), .Z(n167) );
  BUF_X1 U295 ( .A(BTB_PC_From_DE[14]), .Z(n170) );
  BUF_X1 U296 ( .A(BTB_PC_From_DE[15]), .Z(n173) );
  BUF_X1 U297 ( .A(BTB_PC_From_DE[16]), .Z(n176) );
  BUF_X1 U298 ( .A(BTB_PC_From_DE[17]), .Z(n179) );
  BUF_X1 U299 ( .A(BTB_PC_From_DE[18]), .Z(n182) );
  BUF_X1 U300 ( .A(BTB_PC_From_DE[19]), .Z(n185) );
  BUF_X1 U301 ( .A(BTB_PC_From_DE[20]), .Z(n188) );
  BUF_X1 U302 ( .A(BTB_PC_From_DE[21]), .Z(n191) );
  BUF_X1 U303 ( .A(BTB_PC_From_DE[22]), .Z(n194) );
  BUF_X1 U304 ( .A(BTB_PC_From_DE[23]), .Z(n197) );
  BUF_X1 U305 ( .A(BTB_PC_From_DE[24]), .Z(n200) );
  BUF_X1 U306 ( .A(BTB_PC_From_DE[25]), .Z(n203) );
  BUF_X1 U307 ( .A(BTB_PC_From_DE[26]), .Z(n206) );
  BUF_X1 U308 ( .A(BTB_PC_From_DE[27]), .Z(n209) );
  BUF_X1 U309 ( .A(BTB_PC_From_DE[28]), .Z(n212) );
  BUF_X1 U310 ( .A(BTB_PC_From_DE[29]), .Z(n215) );
  BUF_X1 U311 ( .A(BTB_target_From_DE[0]), .Z(n32) );
  BUF_X1 U312 ( .A(n5), .Z(n11) );
  BUF_X1 U313 ( .A(n5), .Z(n12) );
  BUF_X1 U314 ( .A(n5), .Z(n13) );
  BUF_X1 U315 ( .A(s_selmuxes_Fencoder_Tmuxes[2]), .Z(n26) );
  BUF_X1 U316 ( .A(n3), .Z(n14) );
  NOR3_X1 U317 ( .A1(n6), .A2(s_HIT_miss_Freg_Txor), .A3(BTB_restore), .ZN(n3)
         );
  INV_X1 U318 ( .A(BTB_is_branch), .ZN(n6) );
  BUF_X1 U319 ( .A(BTB_rst), .Z(n326) );
  BUF_X1 U320 ( .A(BTB_rst), .Z(n327) );
  BUF_X1 U321 ( .A(BTB_rst), .Z(n325) );
  CLKBUF_X1 U322 ( .A(s_selmuxes_Fencoder_Tmuxes[1]), .Z(n23) );
  CLKBUF_X1 U323 ( .A(s_selmuxes_Fencoder_Tmuxes[1]), .Z(n24) );
  CLKBUF_X1 U324 ( .A(s_selmuxes_Fencoder_Tmuxes[1]), .Z(n25) );
  INV_X1 U325 ( .A(n324), .ZN(n318) );
  INV_X1 U326 ( .A(n324), .ZN(n319) );
  INV_X1 U327 ( .A(n324), .ZN(n320) );
  INV_X1 U328 ( .A(n324), .ZN(n321) );
  INV_X1 U329 ( .A(n324), .ZN(n322) );
  INV_X1 U330 ( .A(n324), .ZN(n323) );
endmodule


module BTB_misprediction_manager_NBIT_PC32 ( BMM_clk, BMM_reset, BMM_enable, 
        BMM_restore, BMM_PC, BMM_NPC, BMM_computed_PC, BMM_is_branch, 
        BMM_branch_taken, BMM_PC_BTB, BMM_NPC_BTB, BMM_computed_PC_BTB, 
        BMM_restore_BTB, BMM_is_branch_BTB, BMM_branch_taken_BTB );
  input [31:0] BMM_PC;
  input [31:0] BMM_NPC;
  input [31:0] BMM_computed_PC;
  output [31:0] BMM_PC_BTB;
  output [31:0] BMM_NPC_BTB;
  output [31:0] BMM_computed_PC_BTB;
  input BMM_clk, BMM_reset, BMM_enable, BMM_restore, BMM_is_branch,
         BMM_branch_taken;
  output BMM_restore_BTB, BMM_is_branch_BTB, BMM_branch_taken_BTB;
  wire   s_restore, s_rst, s_cnt_out_xored, s_not_cnt_out_xored,
         s_restore_Freg_Tmux, s_is_branch_Freg_Tmux, s_branch_taken_Freg_Tmux,
         s_not_branch_taken;
  wire   [1:0] s_cnt_out;
  wire   [31:0] s_pc_Freg_Tmux;
  wire   [31:0] s_npc_Freg_Tmux;
  wire   [31:0] s_computed_pc_Freg_Tmux;

  Reg1Bit_14 RESTORE_REG ( .clk(BMM_clk), .reset(BMM_reset), .data_in(
        BMM_restore), .enable(BMM_enable), .load(1'b1), .data_out(s_restore)
         );
  SAT_Counter_N2 CNT ( .SAT_clk(BMM_clk), .SAT_reset(BMM_reset), .SAT_enable(
        BMM_enable), .SAT_Ud(1'b0), .SAT_update(1'b1), .SAT_setToDef(s_rst), 
        .SAT_SO(s_cnt_out) );
  NRegister_N32_110 REG_PC ( .clk(BMM_clk), .reset(BMM_reset), .data_in(BMM_PC), .enable(s_not_cnt_out_xored), .load(1'b1), .data_out(s_pc_Freg_Tmux) );
  NRegister_N32_109 REG_NPC ( .clk(BMM_clk), .reset(BMM_reset), .data_in(
        BMM_NPC), .enable(s_not_cnt_out_xored), .load(1'b1), .data_out(
        s_npc_Freg_Tmux) );
  NRegister_N32_108 REG_computed_PC ( .clk(BMM_clk), .reset(BMM_reset), 
        .data_in(BMM_computed_PC), .enable(s_not_cnt_out_xored), .load(1'b1), 
        .data_out(s_computed_pc_Freg_Tmux) );
  Reg1Bit_13 REG_RESTORE ( .clk(BMM_clk), .reset(BMM_reset), .data_in(
        BMM_restore), .enable(s_not_cnt_out_xored), .load(1'b1), .data_out(
        s_restore_Freg_Tmux) );
  Reg1Bit_12 IS_BRANCH_REG ( .clk(BMM_clk), .reset(BMM_reset), .data_in(
        BMM_is_branch), .enable(s_not_cnt_out_xored), .load(1'b1), .data_out(
        s_is_branch_Freg_Tmux) );
  Reg1Bit_11 BRANCH_TAKEN_REG ( .clk(BMM_clk), .reset(BMM_reset), .data_in(
        BMM_branch_taken), .enable(s_not_cnt_out_xored), .load(1'b1), 
        .data_out(s_branch_taken_Freg_Tmux) );
  Mux_NBit_2x1_NBIT_IN32_127 MUX_PC ( .port0(BMM_PC), .port1(s_npc_Freg_Tmux), 
        .sel(s_cnt_out_xored), .portY(BMM_PC_BTB) );
  Mux_NBit_2x1_NBIT_IN32_126 MUX_NPC ( .port0(BMM_NPC), .port1(s_pc_Freg_Tmux), 
        .sel(s_cnt_out_xored), .portY(BMM_NPC_BTB) );
  Mux_NBit_2x1_NBIT_IN32_125 MUX_computed_PC ( .port0(BMM_computed_PC), 
        .port1(s_computed_pc_Freg_Tmux), .sel(s_cnt_out_xored), .portY(
        BMM_computed_PC_BTB) );
  Mux_1Bit_2X1_0 MUX_RESTORE ( .port0(s_restore), .port1(s_restore_Freg_Tmux), 
        .sel(s_cnt_out_xored), .portY(BMM_restore_BTB) );
  Mux_1Bit_2X1_7 MUX_IS_BRANCH ( .port0(BMM_is_branch), .port1(
        s_is_branch_Freg_Tmux), .sel(s_cnt_out_xored), .portY(
        BMM_is_branch_BTB) );
  Mux_1Bit_2X1_6 MUX_BRANCH_TAKEN ( .port0(BMM_branch_taken), .port1(
        s_not_branch_taken), .sel(s_cnt_out_xored), .portY(
        BMM_branch_taken_BTB) );
  INV_X1 U3 ( .A(s_not_cnt_out_xored), .ZN(s_cnt_out_xored) );
  INV_X1 U4 ( .A(s_branch_taken_Freg_Tmux), .ZN(s_not_branch_taken) );
  XNOR2_X1 U5 ( .A(s_cnt_out[1]), .B(s_cnt_out[0]), .ZN(s_not_cnt_out_xored)
         );
  OR2_X1 U6 ( .A1(BMM_reset), .A2(s_restore), .ZN(s_rst) );
endmodule


module NRegister_N32_0 ( clk, reset, data_in, enable, load, data_out );
  input [31:0] data_in;
  output [31:0] data_out;
  input clk, reset, enable, load;
  wire   n68, n69, n70, n71, n72, n73, n74, n75, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n85, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95,
         n96, n97, n98, n100, net106709, net106710, net106711, net106712,
         net106713, net106714, net106715, net106716, net106717, net106718,
         net106719, net106720, net106721, net106722, net106723, net106724,
         net106725, net106726, net106727, net106728, net106729, net106730,
         net106731, net106732, net106733, net106734, net106735, net106736,
         net106737, net106738, net106739, net106740, n35, n36, n38, n39, n40,
         n41, n42, n43, n44, n45, n46, n47, n48, n49, n50, n51, n52, n53, n54,
         n55, n56, n57, n58, n59, n60, n61, n62, n63, n64, n65, n66, n67, n101,
         n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14;

  DFFR_X1 \data_out_reg[31]  ( .D(n100), .CK(clk), .RN(n13), .Q(data_out[31]), 
        .QN(net106740) );
  DFFR_X1 \data_out_reg[30]  ( .D(n98), .CK(clk), .RN(n13), .Q(data_out[30]), 
        .QN(net106739) );
  DFFR_X1 \data_out_reg[29]  ( .D(n97), .CK(clk), .RN(n11), .Q(data_out[29]), 
        .QN(net106738) );
  DFFR_X1 \data_out_reg[28]  ( .D(n96), .CK(clk), .RN(n11), .Q(data_out[28]), 
        .QN(net106737) );
  DFFR_X1 \data_out_reg[27]  ( .D(n95), .CK(clk), .RN(n11), .Q(data_out[27]), 
        .QN(net106736) );
  DFFR_X1 \data_out_reg[26]  ( .D(n94), .CK(clk), .RN(n11), .Q(data_out[26]), 
        .QN(net106735) );
  DFFR_X1 \data_out_reg[25]  ( .D(n93), .CK(clk), .RN(n11), .Q(data_out[25]), 
        .QN(net106734) );
  DFFR_X1 \data_out_reg[24]  ( .D(n92), .CK(clk), .RN(n13), .Q(data_out[24]), 
        .QN(net106733) );
  DFFR_X1 \data_out_reg[23]  ( .D(n91), .CK(clk), .RN(n11), .Q(data_out[23]), 
        .QN(net106732) );
  DFFR_X1 \data_out_reg[22]  ( .D(n90), .CK(clk), .RN(n11), .Q(data_out[22]), 
        .QN(net106731) );
  DFFR_X1 \data_out_reg[21]  ( .D(n89), .CK(clk), .RN(n11), .Q(data_out[21]), 
        .QN(net106730) );
  DFFR_X1 \data_out_reg[20]  ( .D(n88), .CK(clk), .RN(n11), .Q(data_out[20]), 
        .QN(net106729) );
  DFFR_X1 \data_out_reg[19]  ( .D(n87), .CK(clk), .RN(n11), .Q(data_out[19]), 
        .QN(net106728) );
  DFFR_X1 \data_out_reg[18]  ( .D(n86), .CK(clk), .RN(n12), .Q(data_out[18]), 
        .QN(net106727) );
  DFFR_X1 \data_out_reg[17]  ( .D(n85), .CK(clk), .RN(n12), .Q(data_out[17]), 
        .QN(net106726) );
  DFFR_X1 \data_out_reg[16]  ( .D(n84), .CK(clk), .RN(n12), .Q(data_out[16]), 
        .QN(net106725) );
  DFFR_X1 \data_out_reg[15]  ( .D(n83), .CK(clk), .RN(n12), .Q(data_out[15]), 
        .QN(net106724) );
  DFFR_X1 \data_out_reg[14]  ( .D(n82), .CK(clk), .RN(n13), .Q(data_out[14]), 
        .QN(net106723) );
  DFFR_X1 \data_out_reg[13]  ( .D(n81), .CK(clk), .RN(n13), .Q(data_out[13]), 
        .QN(net106722) );
  DFFR_X1 \data_out_reg[12]  ( .D(n80), .CK(clk), .RN(n12), .Q(data_out[12]), 
        .QN(net106721) );
  DFFR_X1 \data_out_reg[11]  ( .D(n79), .CK(clk), .RN(n12), .Q(data_out[11]), 
        .QN(net106720) );
  DFFR_X1 \data_out_reg[10]  ( .D(n78), .CK(clk), .RN(n11), .Q(data_out[10]), 
        .QN(net106719) );
  DFFR_X1 \data_out_reg[9]  ( .D(n77), .CK(clk), .RN(n13), .Q(data_out[9]), 
        .QN(net106718) );
  DFFR_X1 \data_out_reg[8]  ( .D(n76), .CK(clk), .RN(n13), .Q(data_out[8]), 
        .QN(net106717) );
  DFFR_X1 \data_out_reg[7]  ( .D(n75), .CK(clk), .RN(n11), .Q(data_out[7]), 
        .QN(net106716) );
  DFFR_X1 \data_out_reg[6]  ( .D(n74), .CK(clk), .RN(n12), .Q(data_out[6]), 
        .QN(net106715) );
  DFFR_X1 \data_out_reg[5]  ( .D(n73), .CK(clk), .RN(n12), .Q(data_out[5]), 
        .QN(net106714) );
  DFFR_X1 \data_out_reg[4]  ( .D(n72), .CK(clk), .RN(n12), .Q(data_out[4]), 
        .QN(net106713) );
  DFFR_X1 \data_out_reg[3]  ( .D(n71), .CK(clk), .RN(n12), .Q(data_out[3]), 
        .QN(net106712) );
  DFFR_X1 \data_out_reg[2]  ( .D(n70), .CK(clk), .RN(n12), .Q(data_out[2]), 
        .QN(net106711) );
  DFFR_X1 \data_out_reg[1]  ( .D(n69), .CK(clk), .RN(n12), .Q(data_out[1]), 
        .QN(net106710) );
  DFFR_X1 \data_out_reg[0]  ( .D(n68), .CK(clk), .RN(n13), .Q(data_out[0]), 
        .QN(net106709) );
  INV_X1 U3 ( .A(n10), .ZN(n3) );
  INV_X1 U4 ( .A(n10), .ZN(n2) );
  BUF_X1 U5 ( .A(n35), .Z(n9) );
  BUF_X1 U6 ( .A(n35), .Z(n8) );
  BUF_X1 U7 ( .A(n35), .Z(n7) );
  BUF_X1 U8 ( .A(n35), .Z(n6) );
  BUF_X1 U9 ( .A(n35), .Z(n5) );
  BUF_X1 U10 ( .A(n35), .Z(n4) );
  BUF_X1 U11 ( .A(n35), .Z(n10) );
  BUF_X1 U12 ( .A(n14), .Z(n12) );
  BUF_X1 U13 ( .A(n14), .Z(n11) );
  BUF_X1 U14 ( .A(n14), .Z(n13) );
  NAND2_X1 U15 ( .A1(load), .A2(enable), .ZN(n35) );
  OAI22_X1 U16 ( .A1(n5), .A2(n44), .B1(net106732), .B2(n3), .ZN(n91) );
  INV_X1 U17 ( .A(data_in[23]), .ZN(n44) );
  OAI22_X1 U18 ( .A1(n5), .A2(n43), .B1(net106733), .B2(n2), .ZN(n92) );
  INV_X1 U19 ( .A(data_in[24]), .ZN(n43) );
  OAI22_X1 U20 ( .A1(n5), .A2(n42), .B1(net106734), .B2(n3), .ZN(n93) );
  INV_X1 U21 ( .A(data_in[25]), .ZN(n42) );
  OAI22_X1 U22 ( .A1(n4), .A2(n41), .B1(net106735), .B2(n2), .ZN(n94) );
  INV_X1 U23 ( .A(data_in[26]), .ZN(n41) );
  OAI22_X1 U24 ( .A1(n4), .A2(n40), .B1(net106736), .B2(n3), .ZN(n95) );
  INV_X1 U25 ( .A(data_in[27]), .ZN(n40) );
  OAI22_X1 U26 ( .A1(n4), .A2(n39), .B1(net106737), .B2(n2), .ZN(n96) );
  INV_X1 U27 ( .A(data_in[28]), .ZN(n39) );
  OAI22_X1 U28 ( .A1(n4), .A2(n38), .B1(net106738), .B2(n3), .ZN(n97) );
  INV_X1 U29 ( .A(data_in[29]), .ZN(n38) );
  OAI22_X1 U30 ( .A1(n4), .A2(n36), .B1(net106739), .B2(n2), .ZN(n98) );
  INV_X1 U31 ( .A(data_in[30]), .ZN(n36) );
  OAI22_X1 U32 ( .A1(n10), .A2(n67), .B1(net106709), .B2(n2), .ZN(n68) );
  INV_X1 U33 ( .A(data_in[0]), .ZN(n67) );
  OAI22_X1 U34 ( .A1(n9), .A2(n66), .B1(net106710), .B2(n2), .ZN(n69) );
  INV_X1 U35 ( .A(data_in[1]), .ZN(n66) );
  OAI22_X1 U36 ( .A1(n9), .A2(n65), .B1(net106711), .B2(n2), .ZN(n70) );
  INV_X1 U37 ( .A(data_in[2]), .ZN(n65) );
  OAI22_X1 U38 ( .A1(n9), .A2(n64), .B1(net106712), .B2(n2), .ZN(n71) );
  INV_X1 U39 ( .A(data_in[3]), .ZN(n64) );
  OAI22_X1 U40 ( .A1(n9), .A2(n63), .B1(net106713), .B2(n2), .ZN(n72) );
  INV_X1 U41 ( .A(data_in[4]), .ZN(n63) );
  OAI22_X1 U42 ( .A1(n9), .A2(n62), .B1(net106714), .B2(n2), .ZN(n73) );
  INV_X1 U43 ( .A(data_in[5]), .ZN(n62) );
  OAI22_X1 U44 ( .A1(n8), .A2(n61), .B1(net106715), .B2(n2), .ZN(n74) );
  INV_X1 U45 ( .A(data_in[6]), .ZN(n61) );
  OAI22_X1 U46 ( .A1(n8), .A2(n60), .B1(net106716), .B2(n2), .ZN(n75) );
  INV_X1 U47 ( .A(data_in[7]), .ZN(n60) );
  OAI22_X1 U48 ( .A1(n8), .A2(n59), .B1(net106717), .B2(n2), .ZN(n76) );
  INV_X1 U49 ( .A(data_in[8]), .ZN(n59) );
  OAI22_X1 U50 ( .A1(n8), .A2(n58), .B1(net106718), .B2(n2), .ZN(n77) );
  INV_X1 U51 ( .A(data_in[9]), .ZN(n58) );
  OAI22_X1 U52 ( .A1(n8), .A2(n57), .B1(net106719), .B2(n2), .ZN(n78) );
  INV_X1 U53 ( .A(data_in[10]), .ZN(n57) );
  OAI22_X1 U54 ( .A1(n7), .A2(n56), .B1(net106720), .B2(n3), .ZN(n79) );
  INV_X1 U55 ( .A(data_in[11]), .ZN(n56) );
  OAI22_X1 U56 ( .A1(n7), .A2(n55), .B1(net106721), .B2(n3), .ZN(n80) );
  INV_X1 U57 ( .A(data_in[12]), .ZN(n55) );
  OAI22_X1 U58 ( .A1(n7), .A2(n54), .B1(net106722), .B2(n3), .ZN(n81) );
  INV_X1 U59 ( .A(data_in[13]), .ZN(n54) );
  OAI22_X1 U60 ( .A1(n7), .A2(n53), .B1(net106723), .B2(n3), .ZN(n82) );
  INV_X1 U61 ( .A(data_in[14]), .ZN(n53) );
  OAI22_X1 U62 ( .A1(n7), .A2(n52), .B1(net106724), .B2(n3), .ZN(n83) );
  INV_X1 U63 ( .A(data_in[15]), .ZN(n52) );
  OAI22_X1 U64 ( .A1(n6), .A2(n51), .B1(net106725), .B2(n3), .ZN(n84) );
  INV_X1 U65 ( .A(data_in[16]), .ZN(n51) );
  OAI22_X1 U66 ( .A1(n6), .A2(n50), .B1(net106726), .B2(n3), .ZN(n85) );
  INV_X1 U67 ( .A(data_in[17]), .ZN(n50) );
  OAI22_X1 U68 ( .A1(n6), .A2(n49), .B1(net106727), .B2(n3), .ZN(n86) );
  INV_X1 U69 ( .A(data_in[18]), .ZN(n49) );
  OAI22_X1 U70 ( .A1(n6), .A2(n48), .B1(net106728), .B2(n3), .ZN(n87) );
  INV_X1 U71 ( .A(data_in[19]), .ZN(n48) );
  OAI22_X1 U72 ( .A1(n6), .A2(n47), .B1(net106729), .B2(n3), .ZN(n88) );
  INV_X1 U73 ( .A(data_in[20]), .ZN(n47) );
  OAI22_X1 U74 ( .A1(n5), .A2(n46), .B1(net106730), .B2(n3), .ZN(n89) );
  INV_X1 U75 ( .A(data_in[21]), .ZN(n46) );
  OAI22_X1 U76 ( .A1(n5), .A2(n45), .B1(net106731), .B2(n3), .ZN(n90) );
  INV_X1 U77 ( .A(data_in[22]), .ZN(n45) );
  OAI22_X1 U78 ( .A1(n10), .A2(n101), .B1(net106740), .B2(n2), .ZN(n100) );
  INV_X1 U79 ( .A(data_in[31]), .ZN(n101) );
  INV_X1 U80 ( .A(reset), .ZN(n14) );
endmodule


module ControlUnit ( CU_instr_opcode, CU_instr_func, CU_enable, CU_reset, 
        CU_clk, CU_flush, CU_bubble, CU_CW_DE, CU_CW_EX, CU_CW_MEM, CU_CW_WB, 
        CU_error );
  input [5:0] CU_instr_opcode;
  input [10:0] CU_instr_func;
  output [1:9] CU_CW_DE;
  output [8:16] CU_CW_EX;
  output [17:22] CU_CW_MEM;
  output [23:26] CU_CW_WB;
  input CU_enable, CU_reset, CU_clk, CU_flush, CU_bubble;
  output CU_error;
  wire   s_insert_nop, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n70, n71, n72, n73, n74, n75, n76, n77,
         n78, n79, n80, n81, n82, n83, n84, n85, n86, n87, n88, n89, n90, n91,
         n92, n93, n94, n95, n96, n97, n98, n99, n100, n101, n102, n103, n104,
         n105, n106, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n118, n119, n120, n121, n122, n123, n124, n125, n126,
         n127, n128, n129, n130, n131, n132, n133, n134, n135, n136, n137,
         n138, n139, n140, n141, n142, n143, n144, n145, n146, n147, n148,
         n149, n150, n151, n152, n153, n154, n155, n156, n157, n158, n159,
         n160, n161, n162, n163, n164, n165, n166, n167, n168, n169, n170,
         n171, n172, n173, n174, n175, n176, n177, n178, n179, n180, n181,
         n182, n183, n184, n185, n186, n187, n188, n189, n190, n191, n192,
         n193, n194, n195, n196, n197, n198, n199, n200, n201, n202, n203,
         n204, n205, n206, n207, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n221, n222, n223, n225, n226,
         n227, n228, n229, n230, n231, n232, n224, n233;
  wire   [1:26] s_control_word;
  wire   [1:26] s_cw_bubble;
  wire   [1:26] s_cw_tmp;
  wire   [10:26] s_cw_Fde_Tex;
  wire   [17:26] s_cw_Fex_Tmem;
  wire   [23:26] s_cw_Fmem_Twb;

  NOR3_X2 U143 ( .A1(CU_instr_opcode[4]), .A2(CU_instr_opcode[5]), .A3(n208), 
        .ZN(n161) );
  NAND3_X1 U219 ( .A1(n79), .A2(n80), .A3(n81), .ZN(s_control_word[6]) );
  NAND3_X1 U220 ( .A1(n101), .A2(n100), .A3(n102), .ZN(s_control_word[1]) );
  NAND3_X1 U221 ( .A1(n132), .A2(n133), .A3(n134), .ZN(n105) );
  NAND3_X1 U222 ( .A1(n156), .A2(n157), .A3(n158), .ZN(n153) );
  NAND3_X1 U223 ( .A1(n145), .A2(n77), .A3(n73), .ZN(n170) );
  NAND3_X1 U224 ( .A1(n87), .A2(n124), .A3(n161), .ZN(n75) );
  NAND3_X1 U225 ( .A1(n116), .A2(n181), .A3(n86), .ZN(n179) );
  NAND3_X1 U226 ( .A1(n104), .A2(n188), .A3(n189), .ZN(n187) );
  NAND3_X1 U227 ( .A1(n136), .A2(n193), .A3(CU_instr_func[1]), .ZN(n192) );
  NAND3_X1 U228 ( .A1(n61), .A2(n196), .A3(n197), .ZN(n140) );
  NAND3_X1 U229 ( .A1(CU_instr_func[1]), .A2(n136), .A3(CU_instr_func[0]), 
        .ZN(n197) );
  NAND3_X1 U230 ( .A1(n198), .A2(n188), .A3(n136), .ZN(n61) );
  NAND3_X1 U231 ( .A1(n149), .A2(CU_instr_opcode[0]), .A3(n147), .ZN(n203) );
  NAND3_X1 U232 ( .A1(n149), .A2(CU_instr_opcode[0]), .A3(n161), .ZN(n204) );
  NAND3_X1 U233 ( .A1(CU_instr_func[5]), .A2(n199), .A3(n135), .ZN(n139) );
  NAND3_X1 U234 ( .A1(n199), .A2(n188), .A3(CU_instr_func[5]), .ZN(n196) );
  NAND3_X1 U235 ( .A1(n86), .A2(n117), .A3(n214), .ZN(n131) );
  Mux_NBit_2x1_NBIT_IN26 BUBBLE_MUX ( .port0({s_control_word[1:19], 
        s_control_word[23], s_control_word[21:26]}), .port1({1'b0, 1'b0, 1'b0, 
        s_cw_bubble[4:7], 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b1, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sel(
        s_insert_nop), .portY(s_cw_tmp) );
  NRegister_N26 DE_CW ( .clk(CU_clk), .reset(CU_reset), .data_in(s_cw_tmp), 
        .enable(n224), .load(1'b1), .data_out({CU_CW_DE, s_cw_Fde_Tex}) );
  NRegister_N19 EX_CW ( .clk(CU_clk), .reset(CU_reset), .data_in({
        CU_CW_DE[8:9], s_cw_Fde_Tex}), .enable(n224), .load(1'b1), .data_out({
        CU_CW_EX, s_cw_Fex_Tmem}) );
  NRegister_N10 MEM_CW ( .clk(CU_clk), .reset(CU_reset), .data_in(
        s_cw_Fex_Tmem), .enable(n224), .load(1'b1), .data_out({CU_CW_MEM, 
        s_cw_Fmem_Twb}) );
  NRegister_N4 WB_CW ( .clk(CU_clk), .reset(CU_reset), .data_in(s_cw_Fmem_Twb), 
        .enable(n224), .load(1'b1), .data_out(CU_CW_WB) );
  NAND2_X2 U25 ( .A1(CU_bubble), .A2(n53), .ZN(s_insert_nop) );
  NOR2_X1 U26 ( .A1(n233), .A2(CU_reset), .ZN(n67) );
  INV_X1 U27 ( .A(n104), .ZN(n62) );
  OAI21_X1 U28 ( .B1(n92), .B2(n62), .A(n93), .ZN(s_control_word[2]) );
  INV_X1 U29 ( .A(n66), .ZN(n56) );
  NOR2_X1 U30 ( .A1(n54), .A2(n55), .ZN(s_cw_bubble[7]) );
  OR2_X1 U31 ( .A1(n54), .A2(s_control_word[6]), .ZN(s_cw_bubble[6]) );
  AOI211_X1 U32 ( .C1(n125), .C2(n126), .A(n120), .B(s_control_word[21]), .ZN(
        n93) );
  NOR2_X1 U33 ( .A1(n116), .A2(n125), .ZN(n145) );
  NOR2_X1 U34 ( .A1(n131), .A2(n58), .ZN(n104) );
  OAI21_X1 U35 ( .B1(n85), .B2(n74), .A(n82), .ZN(n66) );
  AOI21_X1 U36 ( .B1(n82), .B2(n83), .A(n58), .ZN(s_control_word[5]) );
  NAND4_X1 U37 ( .A1(n81), .A2(n79), .A3(n111), .A4(n74), .ZN(
        s_control_word[19]) );
  NOR2_X1 U38 ( .A1(n95), .A2(n98), .ZN(s_control_word[26]) );
  NOR2_X1 U39 ( .A1(n128), .A2(n77), .ZN(s_control_word[22]) );
  INV_X1 U40 ( .A(n69), .ZN(n80) );
  INV_X1 U41 ( .A(n148), .ZN(n122) );
  INV_X1 U42 ( .A(n74), .ZN(n86) );
  OAI21_X1 U43 ( .B1(n89), .B2(n58), .A(n93), .ZN(s_control_word[16]) );
  INV_X1 U44 ( .A(n162), .ZN(n109) );
  OAI21_X1 U45 ( .B1(n73), .B2(n95), .A(n97), .ZN(s_control_word[24]) );
  INV_X1 U46 ( .A(s_control_word[26]), .ZN(n97) );
  INV_X1 U47 ( .A(n101), .ZN(n120) );
  NAND2_X1 U48 ( .A1(n147), .A2(n125), .ZN(n82) );
  INV_X1 U49 ( .A(n81), .ZN(n106) );
  INV_X1 U50 ( .A(n150), .ZN(n147) );
  INV_X1 U51 ( .A(n125), .ZN(n85) );
  INV_X1 U52 ( .A(n131), .ZN(n193) );
  INV_X1 U53 ( .A(n83), .ZN(n107) );
  INV_X1 U54 ( .A(n105), .ZN(n92) );
  INV_X1 U55 ( .A(n128), .ZN(n126) );
  INV_X1 U56 ( .A(n100), .ZN(s_control_word[23]) );
  INV_X1 U57 ( .A(n127), .ZN(s_control_word[21]) );
  AOI21_X1 U58 ( .B1(n116), .B2(n126), .A(s_control_word[22]), .ZN(n127) );
  INV_X1 U59 ( .A(n55), .ZN(s_control_word[7]) );
  INV_X1 U60 ( .A(n189), .ZN(n157) );
  INV_X1 U61 ( .A(n210), .ZN(n225) );
  INV_X1 U62 ( .A(n53), .ZN(n54) );
  AND2_X1 U63 ( .A1(n53), .A2(s_control_word[5]), .ZN(s_cw_bubble[5]) );
  AND2_X1 U64 ( .A1(n53), .A2(s_control_word[4]), .ZN(s_cw_bubble[4]) );
  NOR4_X1 U65 ( .A1(n141), .A2(n142), .A3(n143), .A4(n144), .ZN(n81) );
  OAI211_X1 U66 ( .C1(n76), .C2(n145), .A(n146), .B(n82), .ZN(n144) );
  AOI22_X1 U67 ( .A1(n87), .A2(n148), .B1(n149), .B2(n63), .ZN(n146) );
  NOR2_X1 U68 ( .A1(n124), .A2(n212), .ZN(n116) );
  NOR2_X1 U69 ( .A1(n72), .A2(n124), .ZN(n125) );
  INV_X1 U70 ( .A(n67), .ZN(n58) );
  NOR3_X1 U71 ( .A1(n121), .A2(n124), .A3(n122), .ZN(n90) );
  NOR3_X1 U72 ( .A1(n208), .A2(n222), .A3(n223), .ZN(n148) );
  NOR2_X1 U73 ( .A1(n162), .A2(n96), .ZN(n73) );
  NOR2_X1 U74 ( .A1(n124), .A2(n178), .ZN(n162) );
  NOR3_X1 U75 ( .A1(n106), .A2(n59), .A3(n130), .ZN(n89) );
  OAI221_X1 U76 ( .B1(n74), .B2(n85), .C1(n131), .C2(n92), .A(n111), .ZN(n130)
         );
  NAND2_X1 U77 ( .A1(n171), .A2(n222), .ZN(n74) );
  OAI221_X1 U78 ( .B1(n165), .B2(n122), .C1(n145), .C2(n166), .A(n75), .ZN(
        n164) );
  NOR2_X1 U79 ( .A1(n125), .A2(n162), .ZN(n165) );
  OAI221_X1 U80 ( .B1(n206), .B2(n58), .C1(n62), .C2(n196), .A(n101), .ZN(
        s_control_word[11]) );
  AOI21_X1 U81 ( .B1(n96), .B2(n161), .A(n191), .ZN(n206) );
  OAI21_X1 U82 ( .B1(n64), .B2(n87), .A(n163), .ZN(n78) );
  NAND4_X1 U83 ( .A1(n210), .A2(n86), .A3(n67), .A4(n116), .ZN(n101) );
  AOI22_X1 U84 ( .A1(n96), .A2(n86), .B1(n87), .B2(n63), .ZN(n83) );
  OAI211_X1 U85 ( .C1(n73), .C2(n122), .A(n176), .B(n75), .ZN(n142) );
  OAI21_X1 U86 ( .B1(n117), .B2(n177), .A(n161), .ZN(n176) );
  OAI22_X1 U87 ( .A1(n60), .A2(n58), .B1(n61), .B2(n62), .ZN(s_control_word[8]) );
  AOI211_X1 U88 ( .C1(n63), .C2(n64), .A(n65), .B(n66), .ZN(n60) );
  AOI21_X1 U89 ( .B1(n205), .B2(n116), .A(n173), .ZN(n110) );
  NOR2_X1 U90 ( .A1(n155), .A2(n185), .ZN(n189) );
  OAI21_X1 U91 ( .B1(n212), .B2(n166), .A(n78), .ZN(n143) );
  OAI21_X1 U92 ( .B1(n198), .B2(n196), .A(n139), .ZN(n182) );
  AOI21_X1 U93 ( .B1(n84), .B2(n56), .A(n58), .ZN(s_control_word[4]) );
  OAI21_X1 U94 ( .B1(n63), .B2(n86), .A(n87), .ZN(n84) );
  XNOR2_X1 U95 ( .A(n181), .B(n155), .ZN(n159) );
  INV_X1 U96 ( .A(n161), .ZN(n76) );
  NOR3_X1 U97 ( .A1(n179), .A2(n155), .A3(n180), .ZN(n174) );
  AOI211_X1 U98 ( .C1(n135), .C2(n136), .A(n137), .B(n138), .ZN(n134) );
  INV_X1 U99 ( .A(n140), .ZN(n133) );
  INV_X1 U100 ( .A(n139), .ZN(n138) );
  NOR2_X1 U101 ( .A1(n180), .A2(n159), .ZN(n210) );
  NOR2_X1 U102 ( .A1(n116), .A2(n117), .ZN(n98) );
  AOI21_X1 U103 ( .B1(n56), .B2(n57), .A(n58), .ZN(s_control_word[9]) );
  INV_X1 U104 ( .A(n59), .ZN(n57) );
  AOI21_X1 U105 ( .B1(n88), .B2(n89), .A(n58), .ZN(s_control_word[3]) );
  NOR2_X1 U106 ( .A1(n90), .A2(n91), .ZN(n88) );
  AOI21_X1 U107 ( .B1(n77), .B2(n94), .A(n95), .ZN(s_control_word[25]) );
  INV_X1 U108 ( .A(n96), .ZN(n94) );
  NAND2_X1 U109 ( .A1(n67), .A2(n99), .ZN(n95) );
  OAI211_X1 U110 ( .C1(n132), .C2(n62), .A(n209), .B(n101), .ZN(
        s_control_word[10]) );
  OAI21_X1 U111 ( .B1(n211), .B2(n143), .A(n67), .ZN(n209) );
  AOI21_X1 U112 ( .B1(n73), .B2(n72), .A(n122), .ZN(n211) );
  NAND2_X1 U113 ( .A1(n67), .A2(n69), .ZN(n100) );
  OAI21_X1 U114 ( .B1(n186), .B2(n58), .A(n187), .ZN(s_control_word[13]) );
  AOI211_X1 U115 ( .C1(n163), .C2(n190), .A(n191), .B(n65), .ZN(n186) );
  INV_X1 U116 ( .A(n166), .ZN(n163) );
  INV_X1 U117 ( .A(n190), .ZN(n212) );
  NAND2_X1 U118 ( .A1(n99), .A2(n170), .ZN(n111) );
  INV_X1 U119 ( .A(n117), .ZN(n77) );
  NAND2_X1 U120 ( .A1(n67), .A2(n68), .ZN(n55) );
  OR4_X1 U121 ( .A1(n69), .A2(n59), .A3(n70), .A4(n71), .ZN(n68) );
  OAI21_X1 U122 ( .B1(n76), .B2(n77), .A(n78), .ZN(n70) );
  AOI22_X1 U123 ( .A1(n72), .A2(n73), .B1(n74), .B2(n75), .ZN(n71) );
  NAND2_X1 U124 ( .A1(n67), .A2(n129), .ZN(n128) );
  NAND2_X1 U125 ( .A1(n114), .A2(n208), .ZN(n150) );
  AOI22_X1 U126 ( .A1(n67), .A2(n103), .B1(n104), .B2(n105), .ZN(n102) );
  OR3_X1 U127 ( .A1(n106), .A2(n107), .A3(n108), .ZN(n103) );
  OAI21_X1 U128 ( .B1(n109), .B2(n74), .A(n110), .ZN(n108) );
  OAI21_X1 U129 ( .B1(n171), .B2(n163), .A(n149), .ZN(n218) );
  INV_X1 U130 ( .A(n87), .ZN(n72) );
  NOR2_X1 U131 ( .A1(n178), .A2(n166), .ZN(n175) );
  INV_X1 U132 ( .A(n183), .ZN(n156) );
  NAND2_X1 U133 ( .A1(n169), .A2(n111), .ZN(n69) );
  OAI21_X1 U134 ( .B1(n117), .B2(n172), .A(n129), .ZN(n169) );
  INV_X1 U135 ( .A(n145), .ZN(n172) );
  INV_X1 U136 ( .A(n121), .ZN(n149) );
  AND2_X1 U137 ( .A1(n199), .A2(n200), .ZN(n136) );
  INV_X1 U138 ( .A(n137), .ZN(n185) );
  AND2_X1 U139 ( .A1(n117), .A2(n205), .ZN(n173) );
  INV_X1 U140 ( .A(n207), .ZN(n191) );
  AOI22_X1 U141 ( .A1(n177), .A2(n161), .B1(n182), .B2(n193), .ZN(n207) );
  INV_X1 U142 ( .A(n178), .ZN(n64) );
  AND2_X1 U144 ( .A1(n112), .A2(n113), .ZN(n79) );
  NOR4_X1 U145 ( .A1(n114), .A2(n90), .A3(n91), .A4(n115), .ZN(n113) );
  NOR4_X1 U146 ( .A1(n59), .A2(n58), .A3(n107), .A4(n118), .ZN(n112) );
  AOI21_X1 U147 ( .B1(n98), .B2(n109), .A(n74), .ZN(n115) );
  INV_X1 U148 ( .A(n119), .ZN(s_control_word[18]) );
  AOI21_X1 U149 ( .B1(n67), .B2(n91), .A(n120), .ZN(n119) );
  INV_X1 U150 ( .A(n123), .ZN(s_control_word[17]) );
  AOI21_X1 U151 ( .B1(n67), .B2(n90), .A(n120), .ZN(n123) );
  NOR2_X1 U152 ( .A1(CU_reset), .A2(CU_flush), .ZN(n53) );
  NOR4_X1 U153 ( .A1(n155), .A2(n200), .A3(n160), .A4(CU_instr_func[1]), .ZN(
        n183) );
  NOR2_X1 U154 ( .A1(n212), .A2(CU_instr_opcode[0]), .ZN(n117) );
  NOR3_X1 U155 ( .A1(n121), .A2(CU_instr_opcode[0]), .A3(n122), .ZN(n91) );
  NOR2_X1 U156 ( .A1(n213), .A2(CU_instr_opcode[2]), .ZN(n87) );
  NOR3_X1 U157 ( .A1(n222), .A2(CU_instr_opcode[4]), .A3(n208), .ZN(n129) );
  NOR2_X1 U158 ( .A1(n178), .A2(CU_instr_opcode[0]), .ZN(n96) );
  NOR3_X1 U159 ( .A1(CU_instr_func[6]), .A2(CU_instr_func[10]), .A3(n232), 
        .ZN(n214) );
  OR3_X1 U160 ( .A1(CU_instr_func[9]), .A2(CU_instr_func[8]), .A3(
        CU_instr_func[7]), .ZN(n232) );
  NOR3_X1 U161 ( .A1(CU_instr_func[2]), .A2(CU_instr_func[4]), .A3(n200), .ZN(
        n137) );
  NOR3_X1 U162 ( .A1(n222), .A2(CU_instr_opcode[3]), .A3(n223), .ZN(n205) );
  NOR2_X1 U163 ( .A1(n150), .A2(CU_instr_opcode[0]), .ZN(n63) );
  NOR3_X1 U164 ( .A1(CU_instr_func[3]), .A2(CU_instr_func[4]), .A3(n160), .ZN(
        n199) );
  OAI221_X1 U165 ( .B1(n167), .B2(n62), .C1(n168), .C2(n58), .A(n100), .ZN(
        s_control_word[14]) );
  NOR3_X1 U166 ( .A1(n182), .A2(n183), .A3(n184), .ZN(n167) );
  NOR4_X1 U167 ( .A1(n173), .A2(n174), .A3(n175), .A4(n142), .ZN(n168) );
  NOR3_X1 U168 ( .A1(n185), .A2(CU_instr_func[3]), .A3(CU_instr_func[0]), .ZN(
        n184) );
  NOR2_X1 U169 ( .A1(CU_instr_opcode[2]), .A2(CU_instr_opcode[1]), .ZN(n190)
         );
  NOR2_X1 U170 ( .A1(n188), .A2(CU_instr_func[0]), .ZN(n135) );
  NOR2_X1 U171 ( .A1(n223), .A2(CU_instr_opcode[5]), .ZN(n114) );
  OAI22_X1 U172 ( .A1(n194), .A2(n58), .B1(n195), .B2(n62), .ZN(
        s_control_word[12]) );
  AOI221_X1 U173 ( .B1(n183), .B2(n181), .C1(n189), .C2(CU_instr_func[1]), .A(
        n140), .ZN(n195) );
  NOR3_X1 U174 ( .A1(n201), .A2(n59), .A3(n141), .ZN(n194) );
  OAI21_X1 U175 ( .B1(n76), .B2(n109), .A(n78), .ZN(n201) );
  OAI22_X1 U176 ( .A1(n151), .A2(n58), .B1(n152), .B2(n62), .ZN(
        s_control_word[15]) );
  AOI21_X1 U177 ( .B1(CU_instr_func[0]), .B2(n153), .A(n154), .ZN(n152) );
  AOI221_X1 U178 ( .B1(n125), .B2(n161), .C1(n162), .C2(n163), .A(n164), .ZN(
        n151) );
  AND3_X1 U179 ( .A1(n135), .A2(n155), .A3(n137), .ZN(n154) );
  INV_X1 U180 ( .A(CU_instr_func[2]), .ZN(n160) );
  NOR2_X1 U181 ( .A1(CU_instr_opcode[3]), .A2(CU_instr_opcode[4]), .ZN(n171)
         );
  OAI21_X1 U182 ( .B1(CU_instr_opcode[0]), .B2(n121), .A(n109), .ZN(n177) );
  NAND2_X1 U183 ( .A1(n202), .A2(n203), .ZN(n141) );
  OAI21_X1 U184 ( .B1(n147), .B2(n161), .A(n96), .ZN(n202) );
  INV_X1 U185 ( .A(CU_instr_opcode[0]), .ZN(n124) );
  NAND2_X1 U186 ( .A1(CU_instr_opcode[1]), .A2(CU_instr_opcode[2]), .ZN(n121)
         );
  NAND2_X1 U187 ( .A1(n110), .A2(n204), .ZN(n59) );
  NAND4_X1 U188 ( .A1(n135), .A2(CU_instr_func[2]), .A3(n214), .A4(n200), .ZN(
        n180) );
  INV_X1 U189 ( .A(CU_instr_func[3]), .ZN(n155) );
  NAND4_X1 U190 ( .A1(n218), .A2(n219), .A3(n220), .A4(n221), .ZN(n118) );
  NAND4_X1 U191 ( .A1(CU_instr_opcode[1]), .A2(CU_instr_opcode[5]), .A3(n124), 
        .A4(n223), .ZN(n219) );
  AOI22_X1 U192 ( .A1(n205), .A2(n212), .B1(n129), .B2(CU_instr_opcode[2]), 
        .ZN(n221) );
  OAI21_X1 U193 ( .B1(n147), .B2(n148), .A(n190), .ZN(n220) );
  NAND2_X1 U194 ( .A1(CU_instr_opcode[2]), .A2(n213), .ZN(n178) );
  NAND2_X1 U195 ( .A1(n114), .A2(CU_instr_opcode[3]), .ZN(n166) );
  INV_X1 U196 ( .A(CU_instr_opcode[4]), .ZN(n223) );
  INV_X1 U197 ( .A(CU_instr_opcode[3]), .ZN(n208) );
  INV_X1 U198 ( .A(CU_instr_opcode[5]), .ZN(n222) );
  INV_X1 U199 ( .A(CU_instr_func[5]), .ZN(n200) );
  INV_X1 U200 ( .A(CU_instr_func[1]), .ZN(n188) );
  NAND4_X1 U201 ( .A1(n159), .A2(CU_instr_func[5]), .A3(CU_instr_func[1]), 
        .A4(n160), .ZN(n158) );
  OAI21_X1 U202 ( .B1(n121), .B2(n150), .A(n192), .ZN(n65) );
  INV_X1 U203 ( .A(CU_instr_func[4]), .ZN(n181) );
  AND2_X1 U204 ( .A1(CU_instr_opcode[5]), .A2(n171), .ZN(n99) );
  AND3_X1 U205 ( .A1(n156), .A2(n157), .A3(n215), .ZN(n132) );
  NAND4_X1 U206 ( .A1(CU_instr_func[3]), .A2(CU_instr_func[5]), .A3(
        CU_instr_func[1]), .A4(n160), .ZN(n215) );
  INV_X1 U207 ( .A(CU_instr_opcode[1]), .ZN(n213) );
  INV_X1 U208 ( .A(CU_instr_func[0]), .ZN(n198) );
  AOI211_X1 U209 ( .C1(CU_instr_func[0]), .C2(n188), .A(n160), .B(
        CU_instr_func[3]), .ZN(n227) );
  OAI211_X1 U210 ( .C1(n216), .C2(n74), .A(n67), .B(n217), .ZN(CU_error) );
  INV_X1 U211 ( .A(n118), .ZN(n217) );
  AOI22_X1 U212 ( .A1(n116), .A2(n225), .B1(n117), .B2(n226), .ZN(n216) );
  OAI211_X1 U213 ( .C1(CU_instr_func[5]), .C2(n227), .A(n214), .B(n228), .ZN(
        n226) );
  AOI22_X1 U214 ( .A1(n229), .A2(CU_instr_func[1]), .B1(CU_instr_func[4]), 
        .B2(n230), .ZN(n228) );
  OAI21_X1 U215 ( .B1(CU_instr_func[2]), .B2(CU_instr_func[1]), .A(
        CU_instr_func[3]), .ZN(n230) );
  NOR2_X1 U216 ( .A1(n231), .A2(n160), .ZN(n229) );
  AOI21_X1 U217 ( .B1(CU_instr_func[0]), .B2(CU_instr_func[5]), .A(
        CU_instr_func[3]), .ZN(n231) );
  INV_X1 U218 ( .A(n233), .ZN(n224) );
  INV_X1 U236 ( .A(CU_enable), .ZN(n233) );
endmodule


module Reg1Bit_0 ( clk, reset, data_in, enable, load, data_out );
  input clk, reset, data_in, enable, load;
  output data_out;
  wire   n7, net106708, n4, n5, n2, n3;

  DFFR_X1 data_out_reg ( .D(n7), .CK(clk), .RN(n3), .Q(data_out), .QN(
        net106708) );
  OAI22_X1 U3 ( .A1(net106708), .A2(n4), .B1(n5), .B2(n2), .ZN(n7) );
  INV_X1 U4 ( .A(n5), .ZN(n4) );
  NAND2_X1 U5 ( .A1(load), .A2(enable), .ZN(n5) );
  INV_X1 U6 ( .A(data_in), .ZN(n2) );
  INV_X1 U7 ( .A(reset), .ZN(n3) );
endmodule


module Datapath_NBIT_DATA32_NBIT_IRAM_ADDR5 ( DP_enable, DP_clk, DP_reset, 
        DP_btb_target_prediction, DP_btb_prediction, DP_IR, DP_Rd1, DP_Rd2, 
        DP_Wr, DP_JMP_branch, DP_sign_extender, DP_save_PC, 
        DP_Shift_Amount_sel, DP_use_immediate, DP_reverse_operands, 
        DP_ALU_Opcode, DP_EX_enable, DP_UUW_sel, DP_Store_reduce, 
        DP_Store_BYTE_half, DP_Load_data_from_DRAM, DP_WB_sel, DP_Load_reduce, 
        DP_Load_BYTE_half, DP_Load_SGN_usg_reduce, DP_insert_bubble, DP_PC, 
        DP_NPC, DP_IF_ID_instr_is_branch, DP_IR_opcode, DP_IR_func, 
        DP_restore_BTB, DP_branch_taken, DP_computed_new_PC, DP_target, 
        DP_data_to_DRAM, DP_address_to_DRAM );
  input [31:0] DP_btb_target_prediction;
  input [31:0] DP_IR;
  input [1:0] DP_JMP_branch;
  input [1:0] DP_sign_extender;
  input [1:0] DP_Shift_Amount_sel;
  input [5:0] DP_ALU_Opcode;
  input [1:0] DP_UUW_sel;
  input [31:0] DP_Load_data_from_DRAM;
  output [31:0] DP_PC;
  output [31:0] DP_NPC;
  output [5:0] DP_IR_opcode;
  output [10:0] DP_IR_func;
  output [31:0] DP_computed_new_PC;
  output [31:0] DP_target;
  output [31:0] DP_data_to_DRAM;
  output [31:0] DP_address_to_DRAM;
  input DP_enable, DP_clk, DP_reset, DP_btb_prediction, DP_Rd1, DP_Rd2, DP_Wr,
         DP_save_PC, DP_use_immediate, DP_reverse_operands, DP_EX_enable,
         DP_Store_reduce, DP_Store_BYTE_half, DP_WB_sel, DP_Load_reduce,
         DP_Load_BYTE_half, DP_Load_SGN_usg_reduce;
  output DP_insert_bubble, DP_IF_ID_instr_is_branch, DP_restore_BTB,
         DP_branch_taken;
  wire   n46, \DP_IR[31] , \DP_IR[30] , \DP_IR[29] , \DP_IR[28] , \DP_IR[27] ,
         \DP_IR[26] , \DP_IR[10] , \DP_IR[9] , \DP_IR[8] , \DP_IR[7] ,
         \DP_IR[6] , \DP_IR[5] , \DP_IR[4] , \DP_IR[3] , \DP_IR[2] ,
         \DP_IR[1] , \DP_IR[0] , s_branch_taken_Fde, s_jmp_or_brnch_Ffcu_Tde,
         s_stall_Fif, s_btb_prediction, s_is_jalr_or_jal, s_flush,
         s_reset_middle_regs_ID_EX, s_stall_Fde, s_reset_middle_regs_EX_MEM,
         s_sel_regA_PC_mux, s_use_immediate, s_id_ex_is_store,
         s_use_immediate_sel, s_ex_enable, s_reset_middle_regs_MEM_WB,
         s_stall_Fex, s_ex_mem_fwd_mux, s_IR_Fmem_31, s_IR_Fmem_30,
         s_IR_Fmem_29, s_IR_Fmem_28, s_IR_Fmem_27, s_IR_Fmem_26, s_fcu_enable,
         n5, n6, n7, n9, n8, n10, n11, n12, n13, n14, n15, n16, n17, n18, n19,
         n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30, n31, n32, n33,
         n34, n35, n36, n37, n38, n39, n40, n41, n42, n44, n45;
  wire   [31:0] s_IR_Fif;
  wire   [31:0] s_PC_Tde;
  wire   [31:0] s_NPC_Tde;
  wire   [31:0] s_result_Fex_Tmem;
  wire   [1:0] s_if_id_sel_fwx_mux;
  wire   [31:0] s_data_Fwb_Tde;
  wire   [31:0] s_regA_Fde_Tex;
  wire   [31:0] s_regB_Fde_Tex;
  wire   [31:0] s_regI_Fde_Tex;
  wire   [31:0] s_PC_Tex;
  wire   [31:0] s_IR_Fde;
  wire   [31:0] s_opA_Fmux_Tfrw_mux;
  wire   [31:0] s_opB_Fmux_Tfrw_mux;
  wire   [1:0] s_id_ex_sel_fwd_top_mux;
  wire   [31:0] s_data_fwd_top_alu1;
  wire   [31:0] s_data_fwd_top_alu2;
  wire   [31:0] s_data_fwd_top_aluY;
  wire   [1:0] s_id_ex_sel_fwd_bot_mux;
  wire   [31:0] s_data_fwd_bot_alu1;
  wire   [31:0] s_data_fwd_bot_alu2;
  wire   [31:0] s_data_fwd_bot_aluY;
  wire   [31:0] s_opA_Fmux_Tex;
  wire   [31:0] s_opB_Fmux_Tex;
  wire   [4:0] s_SA_Fmux_Tmux1;
  wire   [4:0] s_SA_Fmux_Tmux2;
  wire   [4:0] s_SA_Fmux_Tex;
  wire   [31:0] s_IR_Fex;
  wire   [31:0] s_dataTBStr_Freg_Tmux;
  wire   [31:0] s_data_TBStr_Fmux_Tex;
  wire   [31:0] s_data_Fmem_Twb;
  wire   [31:0] s_bypass_data_Freg_Twb;
  wire   [20:11] s_IR_Fmem;
  wire   SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15;
  assign DP_IR_opcode[5] = \DP_IR[31] ;
  assign \DP_IR[31]  = DP_IR[31];
  assign DP_IR_opcode[4] = \DP_IR[30] ;
  assign \DP_IR[30]  = DP_IR[30];
  assign DP_IR_opcode[3] = \DP_IR[29] ;
  assign \DP_IR[29]  = DP_IR[29];
  assign DP_IR_opcode[2] = \DP_IR[28] ;
  assign \DP_IR[28]  = DP_IR[28];
  assign DP_IR_opcode[1] = \DP_IR[27] ;
  assign \DP_IR[27]  = DP_IR[27];
  assign DP_IR_opcode[0] = \DP_IR[26] ;
  assign \DP_IR[26]  = DP_IR[26];
  assign DP_IR_func[10] = \DP_IR[10] ;
  assign \DP_IR[10]  = DP_IR[10];
  assign DP_IR_func[9] = \DP_IR[9] ;
  assign \DP_IR[9]  = DP_IR[9];
  assign DP_IR_func[8] = \DP_IR[8] ;
  assign \DP_IR[8]  = DP_IR[8];
  assign DP_IR_func[7] = \DP_IR[7] ;
  assign \DP_IR[7]  = DP_IR[7];
  assign DP_IR_func[6] = \DP_IR[6] ;
  assign \DP_IR[6]  = DP_IR[6];
  assign DP_IR_func[5] = \DP_IR[5] ;
  assign \DP_IR[5]  = DP_IR[5];
  assign DP_IR_func[4] = \DP_IR[4] ;
  assign \DP_IR[4]  = DP_IR[4];
  assign DP_IR_func[3] = \DP_IR[3] ;
  assign \DP_IR[3]  = DP_IR[3];
  assign DP_IR_func[2] = \DP_IR[2] ;
  assign \DP_IR[2]  = DP_IR[2];
  assign DP_IR_func[1] = \DP_IR[1] ;
  assign \DP_IR[1]  = DP_IR[1];
  assign DP_IR_func[0] = \DP_IR[0] ;
  assign \DP_IR[0]  = DP_IR[0];

  Fetch_NBIT_PC32_NBIT_IR32 IF_Stage ( .FE_clk(DP_clk), .FE_rst(n44), 
        .FE_enable(DP_enable), .FE_PC_enable(DP_insert_bubble), .FE_PC_clear(
        n44), .FE_IR_enable(DP_insert_bubble), .FE_IR_clear(n44), 
        .FE_btb_target_prediction(DP_btb_target_prediction), 
        .FE_btb_prediction(DP_btb_prediction), .FE_branch_taken(
        s_branch_taken_Fde), .FE_next_instr_is_branch(DP_IF_ID_instr_is_branch), .FE_next_instr_is_jump(s_jmp_or_brnch_Ffcu_Tde), .FE_new_PC_from_DE(
        DP_computed_new_PC), .FE_IR_in({\DP_IR[31] , \DP_IR[30] , \DP_IR[29] , 
        \DP_IR[28] , \DP_IR[27] , \DP_IR[26] , DP_IR[25:11], \DP_IR[10] , 
        \DP_IR[9] , \DP_IR[8] , \DP_IR[7] , \DP_IR[6] , \DP_IR[5] , \DP_IR[4] , 
        \DP_IR[3] , \DP_IR[2] , \DP_IR[1] , \DP_IR[0] }), .FE_restore_BTB(
        DP_restore_BTB), .FE_IR_out(s_IR_Fif), .FE_PC(DP_PC), .FE_NPC(DP_NPC)
         );
  NRegister_N32_118 PC_IF_ID_REG ( .clk(DP_clk), .reset(n44), .data_in(DP_PC), 
        .enable(DP_insert_bubble), .load(1'b1), .data_out(s_PC_Tde) );
  NRegister_N32_117 NPC_IF_ID_REG ( .clk(DP_clk), .reset(n44), .data_in(DP_NPC), .enable(DP_insert_bubble), .load(1'b1), .data_out(s_NPC_Tde) );
  Reg1Bit_23 stall_IF_ID_REG ( .clk(DP_clk), .reset(n44), .data_in(
        DP_insert_bubble), .enable(DP_enable), .load(1'b1), .data_out(
        s_stall_Fif) );
  Reg1Bit_22 BTB_prediction_IF_ID ( .clk(DP_clk), .reset(n44), .data_in(
        DP_btb_prediction), .enable(DP_enable), .load(1'b1), .data_out(
        s_btb_prediction) );
  Decode_NBIT_PC32_NBIT_IR32_NBIT_ADDR5_NBIT_DATA32 DE_Stage ( .DE_clk(DP_clk), 
        .DE_reset(n44), .DE_enable(DP_enable), .DE_stall(DP_insert_bubble), 
        .DE_IR(s_IR_Fif), .DE_PC(s_PC_Tde), .DE_NPC(s_NPC_Tde), .DE_rd1(DP_Rd1), .DE_rd2(DP_Rd2), .DE_wr(DP_Wr), .DE_data_fex(s_result_Fex_Tmem), 
        .DE_sel_data_forward(s_if_id_sel_fwx_mux), .DE_data_Fwb({n36, n22, n31, 
        n37, n17, n15, s_data_Fwb_Tde[25:23], n10, s_data_Fwb_Tde[21:2], n32, 
        n23}), .DE_signext(DP_sign_extender), .DE_JMP_branch(DP_JMP_branch), 
        .DE_jmp_or_branch(s_jmp_or_brnch_Ffcu_Tde), .DE_save_PC(DP_save_PC), 
        .DE_branch_taken(s_branch_taken_Fde), .DE_new_PC(DP_computed_new_PC), 
        .DE_imm_address(DP_target), .DE_RegA(s_regA_Fde_Tex), .DE_RegB(
        s_regB_Fde_Tex), .DE_RegI(s_regI_Fde_Tex) );
  Reg1Bit_21 flush_ID_EX_REG ( .clk(DP_clk), .reset(n44), .data_in(s_flush), 
        .enable(s_stall_Fif), .load(1'b1), .data_out(s_reset_middle_regs_ID_EX) );
  Reg1Bit_20 stall_ID_EX_REG ( .clk(DP_clk), .reset(n44), .data_in(s_stall_Fif), .enable(DP_enable), .load(1'b1), .data_out(s_stall_Fde) );
  NRegister_N32_116 PC_ID_EX_REG ( .clk(DP_clk), .reset(n44), .data_in(
        s_PC_Tde), .enable(s_stall_Fif), .load(1'b1), .data_out(s_PC_Tex) );
  NRegister_N32_115 IR_ID_EX_REG ( .clk(DP_clk), .reset(
        s_reset_middle_regs_ID_EX), .data_in(s_IR_Fif), .enable(s_stall_Fif), 
        .load(1'b1), .data_out(s_IR_Fde) );
  Reg1Bit_19 RST_ID_EX_REG ( .clk(DP_clk), .reset(n44), .data_in(
        s_reset_middle_regs_ID_EX), .enable(s_stall_Fif), .load(1'b1), 
        .data_out(s_reset_middle_regs_EX_MEM) );
  Mux_NBit_2x1_NBIT_IN32_0 RegA_PC_MUX ( .port0(s_regA_Fde_Tex), .port1(
        s_PC_Tex), .sel(s_sel_regA_PC_mux), .portY(s_opA_Fmux_Tfrw_mux) );
  Reg1Bit_18 REGB_IMM_SEL_REG ( .clk(DP_clk), .reset(n44), .data_in(
        DP_use_immediate), .enable(s_stall_Fif), .load(1'b1), .data_out(
        s_use_immediate) );
  Mux_NBit_2x1_NBIT_IN32_137 RegB_Imm_MUX ( .port0(s_regB_Fde_Tex), .port1(
        s_regI_Fde_Tex), .sel(s_use_immediate_sel), .portY(s_opB_Fmux_Tfrw_mux) );
  Mux_NBit_2x1_NBIT_IN32_136 REG_EX_MEM_TOP_MUX ( .port0(s_opA_Fmux_Tfrw_mux), 
        .port1(s_result_Fex_Tmem), .sel(s_id_ex_sel_fwd_top_mux[0]), .portY(
        s_data_fwd_top_alu1) );
  Mux_NBit_2x1_NBIT_IN32_135 MEM_WB_NULL_TOP_MUX ( .port0(s_data_Fwb_Tde), 
        .port1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sel(
        s_id_ex_sel_fwd_top_mux[0]), .portY(s_data_fwd_top_alu2) );
  Mux_NBit_2x1_NBIT_IN32_134 FWD_TOP_MUX ( .port0(s_data_fwd_top_alu1), 
        .port1(s_data_fwd_top_alu2), .sel(s_id_ex_sel_fwd_top_mux[1]), .portY(
        s_data_fwd_top_aluY) );
  Mux_NBit_2x1_NBIT_IN32_133 REG_EX_MEM_BOT_MUX ( .port0(s_opB_Fmux_Tfrw_mux), 
        .port1(s_result_Fex_Tmem), .sel(s_id_ex_sel_fwd_bot_mux[0]), .portY(
        s_data_fwd_bot_alu1) );
  Mux_NBit_2x1_NBIT_IN32_132 MEM_WB_NULL_BOT_MUX ( .port0(s_data_Fwb_Tde), 
        .port1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sel(
        s_id_ex_sel_fwd_bot_mux[0]), .portY(s_data_fwd_bot_alu2) );
  Mux_NBit_2x1_NBIT_IN32_131 FWD_BOT_MUX ( .port0(s_data_fwd_bot_alu1), 
        .port1(s_data_fwd_bot_alu2), .sel(s_id_ex_sel_fwd_bot_mux[1]), .portY(
        s_data_fwd_bot_aluY) );
  Mux_NBit_2x1_NBIT_IN32_130 REVERSE_TOP_MUX ( .port0({s_data_fwd_top_aluY[31], 
        n16, n30, n35, s_data_fwd_top_aluY[27:0]}), .port1({n8, n28, n26, 
        s_data_fwd_bot_aluY[28], n11, s_data_fwd_bot_aluY[26:0]}), .sel(
        DP_reverse_operands), .portY(s_opA_Fmux_Tex) );
  Mux_NBit_2x1_NBIT_IN32_129 REVERSE_BOT_MUX ( .port0({
        s_data_fwd_bot_aluY[31:3], n18, n25, n33}), .port1({
        s_data_fwd_top_aluY[31:2], n29, s_data_fwd_top_aluY[0]}), .sel(
        DP_reverse_operands), .portY(s_opB_Fmux_Tex) );
  Mux_NBit_2x1_NBIT_IN5_0 SHIFT_AMOUNT_MUX1 ( .port0({1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0}), .port1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sel(
        DP_Shift_Amount_sel[0]), .portY(s_SA_Fmux_Tmux1) );
  Mux_NBit_2x1_NBIT_IN5_4 SHIFT_AMOUNT_MUX2 ( .port0({s_data_fwd_bot_aluY[4:3], 
        n18, n25, n33}), .port1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .sel(
        DP_Shift_Amount_sel[0]), .portY(s_SA_Fmux_Tmux2) );
  Mux_NBit_2x1_NBIT_IN5_3 SHIFT_AMOUNT_MUX3 ( .port0(s_SA_Fmux_Tmux1), .port1(
        s_SA_Fmux_Tmux2), .sel(DP_Shift_Amount_sel[1]), .portY(s_SA_Fmux_Tex)
         );
  Execute_Stage_NBIT_DATA32_NBIT_BS_AMOUNT5 EX_Stage ( .EX_clk(DP_clk), 
        .EX_reset(s_reset_middle_regs_EX_MEM), .EX_enable(s_ex_enable), 
        .EX_OpA(s_opA_Fmux_Tex), .EX_OpB(s_opB_Fmux_Tex), .EX_Opcode(
        DP_ALU_Opcode), .EX_ShiftAmount(s_SA_Fmux_Tex), .EX_sel_mux_out(
        DP_UUW_sel), .EX_data_out(s_result_Fex_Tmem) );
  Reg1Bit_17 RST_EX_MEM_REG ( .clk(DP_clk), .reset(n44), .data_in(
        s_reset_middle_regs_EX_MEM), .enable(s_stall_Fif), .load(1'b1), 
        .data_out(s_reset_middle_regs_MEM_WB) );
  Reg1Bit_16 stall_EX_MEM_REG ( .clk(DP_clk), .reset(
        s_reset_middle_regs_EX_MEM), .data_in(s_stall_Fde), .enable(DP_enable), 
        .load(1'b1), .data_out(s_stall_Fex) );
  NRegister_N32_114 IR_EX_MEM_REG ( .clk(DP_clk), .reset(
        s_reset_middle_regs_EX_MEM), .data_in({s_IR_Fde[31:26], n19, 
        s_IR_Fde[24], n21, s_IR_Fde[22:21], n14, s_IR_Fde[19:0]}), .enable(
        s_stall_Fde), .load(1'b1), .data_out(s_IR_Fex) );
  NRegister_N32_113 OPB_TO_DRAM_REG ( .clk(DP_clk), .reset(
        s_reset_middle_regs_EX_MEM), .data_in(s_regB_Fde_Tex), .enable(
        s_stall_Fde), .load(1'b1), .data_out(s_dataTBStr_Freg_Tmux) );
  Mux_NBit_2x1_NBIT_IN32_128 DATA_TB_STORED_MUX ( .port0(s_dataTBStr_Freg_Tmux), .port1({n36, n22, n31, n37, n17, n15, s_data_Fwb_Tde[25:23], n10, 
        s_data_Fwb_Tde[21:3], n13, n32, n23}), .sel(s_ex_mem_fwd_mux), .portY(
        s_data_TBStr_Fmux_Tex) );
  Memory_Stage_NBIT_DATA32_NBIT_ADDRESS32 MEM_Stage ( .ME_data_in(
        s_data_TBStr_Fmux_Tex), .ME_address(s_result_Fex_Tmem), .ME_clk(DP_clk), .ME_rst(s_reset_middle_regs_MEM_WB), .ME_enable(DP_enable), .ME_reduce(
        DP_Store_reduce), .ME_BYTE_half(DP_Store_BYTE_half), .ME_data_to_mem(
        DP_data_to_DRAM), .ME_address_to_mem(DP_address_to_DRAM), 
        .ME_data_from_mem(DP_Load_data_from_DRAM), .ME_data_rd_out(
        s_data_Fmem_Twb) );
  Reg1Bit_15 stall_MEM_WB_REG ( .clk(DP_clk), .reset(
        s_reset_middle_regs_MEM_WB), .data_in(s_stall_Fex), .enable(DP_enable), 
        .load(1'b1) );
  NRegister_N32_112 DATA_BYPASS_REG ( .clk(DP_clk), .reset(
        s_reset_middle_regs_MEM_WB), .data_in(s_result_Fex_Tmem), .enable(
        s_stall_Fex), .load(1'b1), .data_out(s_bypass_data_Freg_Twb) );
  NRegister_N32_111 IR_MEM_WB_REG ( .clk(DP_clk), .reset(
        s_reset_middle_regs_MEM_WB), .data_in({s_IR_Fex[31:21], n34, 
        s_IR_Fex[19], n39, n41, n20, n24, n12, n27, n42, n40, s_IR_Fex[10:0]}), 
        .enable(s_stall_Fex), .load(1'b1), .data_out({s_IR_Fmem_31, 
        s_IR_Fmem_30, s_IR_Fmem_29, s_IR_Fmem_28, s_IR_Fmem_27, s_IR_Fmem_26, 
        SYNOPSYS_UNCONNECTED__0, SYNOPSYS_UNCONNECTED__1, 
        SYNOPSYS_UNCONNECTED__2, SYNOPSYS_UNCONNECTED__3, 
        SYNOPSYS_UNCONNECTED__4, s_IR_Fmem, SYNOPSYS_UNCONNECTED__5, 
        SYNOPSYS_UNCONNECTED__6, SYNOPSYS_UNCONNECTED__7, 
        SYNOPSYS_UNCONNECTED__8, SYNOPSYS_UNCONNECTED__9, 
        SYNOPSYS_UNCONNECTED__10, SYNOPSYS_UNCONNECTED__11, 
        SYNOPSYS_UNCONNECTED__12, SYNOPSYS_UNCONNECTED__13, 
        SYNOPSYS_UNCONNECTED__14, SYNOPSYS_UNCONNECTED__15}) );
  WriteBack_Stage_NBIT_DATA32 WB_Stage ( .WB_OpA(s_bypass_data_Freg_Twb), 
        .WB_OpB(s_data_Fmem_Twb), .WB_sel(DP_WB_sel), .WB_reduce(
        DP_Load_reduce), .WB_BYTE_half(DP_Load_BYTE_half), .WB_SGN_usg(
        DP_Load_SGN_usg_reduce), .WB_out(s_data_Fwb_Tde) );
  FCU FRW_CU ( .FCU_enable(s_fcu_enable), .FCU_IF_ID_Op(s_IR_Fif[31:26]), 
        .FCU_ID_EX_Op(s_IR_Fde[31:26]), .FCU_EX_MEM_Op(s_IR_Fex[31:26]), 
        .FCU_MEM_WB_Op({s_IR_Fmem_31, s_IR_Fmem_30, s_IR_Fmem_29, s_IR_Fmem_28, 
        s_IR_Fmem_27, s_IR_Fmem_26}), .FCU_IF_ID_6_10(s_IR_Fif[25:21]), 
        .FCU_IF_ID_11_15(s_IR_Fif[20:16]), .FCU_ID_EX_6_10(s_IR_Fde[25:21]), 
        .FCU_ID_EX_11_15(s_IR_Fde[20:16]), .FCU_ID_EX_16_20(s_IR_Fde[15:11]), 
        .FCU_EX_MEM_11_15(s_IR_Fex[20:16]), .FCU_EX_MEM_16_20(s_IR_Fex[15:11]), 
        .FCU_MEM_WB_11_15(s_IR_Fmem[20:16]), .FCU_MEM_WB_16_20(
        s_IR_Fmem[15:11]), .FCU_IF_ID_MUX(s_if_id_sel_fwx_mux), 
        .FCU_ID_EX_TOP_MUX(s_id_ex_sel_fwd_top_mux), .FCU_ID_EX_BOT_MUX(
        s_id_ex_sel_fwd_bot_mux), .FCU_EX_MEM_MUX(s_ex_mem_fwd_mux), 
        .FCU_IF_ID_is_branch(DP_IF_ID_instr_is_branch), .FCU_ID_EX_is_store(
        s_id_ex_is_store), .FCU_IF_ID_is_branch_or_jmp(s_jmp_or_brnch_Ffcu_Tde), .FCU_IF_ID_is_jmp_r(s_is_jalr_or_jal), .FCU_insert_stall(n46) );
  BUF_X1 U3 ( .A(s_data_fwd_bot_aluY[31]), .Z(n8) );
  AND2_X2 U4 ( .A1(n38), .A2(DP_enable), .ZN(s_fcu_enable) );
  CLKBUF_X1 U5 ( .A(s_data_Fwb_Tde[22]), .Z(n10) );
  CLKBUF_X1 U6 ( .A(s_data_fwd_bot_aluY[27]), .Z(n11) );
  CLKBUF_X1 U7 ( .A(s_IR_Fex[14]), .Z(n12) );
  CLKBUF_X1 U8 ( .A(s_data_Fwb_Tde[2]), .Z(n13) );
  CLKBUF_X1 U9 ( .A(s_IR_Fde[20]), .Z(n14) );
  CLKBUF_X1 U10 ( .A(s_data_Fwb_Tde[26]), .Z(n15) );
  CLKBUF_X1 U11 ( .A(s_data_fwd_top_aluY[30]), .Z(n16) );
  CLKBUF_X1 U12 ( .A(s_data_Fwb_Tde[27]), .Z(n17) );
  CLKBUF_X1 U13 ( .A(s_data_fwd_bot_aluY[2]), .Z(n18) );
  CLKBUF_X1 U14 ( .A(s_IR_Fde[25]), .Z(n19) );
  CLKBUF_X1 U15 ( .A(s_IR_Fex[16]), .Z(n20) );
  CLKBUF_X1 U16 ( .A(s_IR_Fde[23]), .Z(n21) );
  CLKBUF_X1 U17 ( .A(s_data_Fwb_Tde[30]), .Z(n22) );
  CLKBUF_X1 U18 ( .A(s_data_Fwb_Tde[0]), .Z(n23) );
  CLKBUF_X1 U19 ( .A(s_IR_Fex[15]), .Z(n24) );
  CLKBUF_X1 U20 ( .A(s_data_fwd_bot_aluY[1]), .Z(n25) );
  CLKBUF_X1 U21 ( .A(s_data_fwd_bot_aluY[29]), .Z(n26) );
  CLKBUF_X1 U22 ( .A(s_IR_Fex[13]), .Z(n27) );
  CLKBUF_X1 U23 ( .A(s_data_fwd_bot_aluY[30]), .Z(n28) );
  CLKBUF_X1 U24 ( .A(s_data_fwd_top_aluY[1]), .Z(n29) );
  CLKBUF_X1 U25 ( .A(s_data_fwd_top_aluY[29]), .Z(n30) );
  CLKBUF_X1 U26 ( .A(s_data_Fwb_Tde[29]), .Z(n31) );
  CLKBUF_X1 U27 ( .A(s_data_Fwb_Tde[1]), .Z(n32) );
  CLKBUF_X1 U28 ( .A(s_data_fwd_bot_aluY[0]), .Z(n33) );
  CLKBUF_X1 U29 ( .A(s_IR_Fex[20]), .Z(n34) );
  CLKBUF_X1 U30 ( .A(s_data_fwd_top_aluY[28]), .Z(n35) );
  CLKBUF_X1 U31 ( .A(s_data_Fwb_Tde[31]), .Z(n36) );
  CLKBUF_X1 U32 ( .A(s_data_Fwb_Tde[28]), .Z(n37) );
  INV_X1 U33 ( .A(DP_reset), .ZN(n38) );
  INV_X1 U34 ( .A(n45), .ZN(n44) );
  INV_X1 U35 ( .A(n6), .ZN(s_sel_regA_PC_mux) );
  BUF_X1 U36 ( .A(n46), .Z(DP_insert_bubble) );
  INV_X1 U37 ( .A(n5), .ZN(s_use_immediate_sel) );
  OAI21_X1 U38 ( .B1(s_id_ex_is_store), .B2(s_use_immediate), .A(n6), .ZN(n5)
         );
  INV_X1 U39 ( .A(DP_reset), .ZN(n45) );
  AND2_X1 U40 ( .A1(DP_EX_enable), .A2(DP_enable), .ZN(s_ex_enable) );
  OAI21_X1 U41 ( .B1(s_is_jalr_or_jal), .B2(n7), .A(n45), .ZN(s_flush) );
  XNOR2_X1 U42 ( .A(s_branch_taken_Fde), .B(s_btb_prediction), .ZN(n7) );
  INV_X1 U43 ( .A(n9), .ZN(DP_branch_taken) );
  OAI21_X1 U44 ( .B1(s_branch_taken_Fde), .B2(s_btb_prediction), .A(
        s_jmp_or_brnch_Ffcu_Tde), .ZN(n9) );
  NAND2_X1 U45 ( .A1(DP_Shift_Amount_sel[1]), .A2(DP_Shift_Amount_sel[0]), 
        .ZN(n6) );
  CLKBUF_X1 U46 ( .A(s_IR_Fex[18]), .Z(n39) );
  CLKBUF_X1 U47 ( .A(s_IR_Fex[11]), .Z(n40) );
  CLKBUF_X1 U48 ( .A(s_IR_Fex[17]), .Z(n41) );
  CLKBUF_X1 U49 ( .A(s_IR_Fex[12]), .Z(n42) );
endmodule


module DLX_Core ( DLX_clk, DLX_reset, DLX_enable, DLX_IR, DLX_read_data, 
        DLX_written_data, DLX_address_written_data, DLX_PC, DLX_enable_DRAM, 
        DLX_RD_wr_DRAM, DLX_error );
  input [31:0] DLX_IR;
  input [31:0] DLX_read_data;
  output [31:0] DLX_written_data;
  output [31:0] DLX_address_written_data;
  output [31:0] DLX_PC;
  input DLX_clk, DLX_reset, DLX_enable;
  output DLX_enable_DRAM, DLX_RD_wr_DRAM, DLX_error;
  wire   s_save_PC_Fcu_Tdp, s_use_immediate_Fcu_Tdp, s_MEM_cw_Fcu_Tdp_21,
         s_MEM_cw_Fcu_Tdp_22, s_insert_bubble_Fdp_Tcu,
         s_IFID_istr_is_brnch_Fdp_Tbmm, s_restore_Fdp_Tbmm,
         s_branch_taken_Fdp_Tdp_cu, s_btb_prediction_Fbtb_Treg,
         s_btb_prediction_Freg_Tcu, s_flush, s_restore_Fbmm_Tbtb,
         s_IFID_istr_is_brnch_Fbmm_Tbtb, s_branch_taken_Fd_bmm_Tbtb, n5, n6,
         n7;
  wire   [1:9] s_DE_cw_Fcu_Tdp;
  wire   [31:0] s_target_prediction_Fbtb_Tdp;
  wire   [8:16] s_EX_cw_Fcu_Tdp;
  wire   [17:18] s_MEM_cw_Fcu_Tdp;
  wire   [23:26] s_WB_cw_Fcu_Tdp;
  wire   [5:0] s_IR_opcode_Fdp_Tcu;
  wire   [10:0] s_IR_func_Fdp_Tcu;
  wire   [31:0] s_computed_NPC_Fdp_Tbmm;
  wire   [31:0] s_NPC_Fdp_Tbmm;
  wire   [31:0] s_PC_Fbmm_Tbtb;
  wire   [31:0] s_NPC_Fbmm_Tbtb;
  wire   [31:0] s_computed_NPC_Fbmm_Tbtb;

  XOR2_X1 U8 ( .A(s_branch_taken_Fdp_Tdp_cu), .B(n5), .Z(s_flush) );
  XOR2_X1 U9 ( .A(s_restore_Fdp_Tbmm), .B(s_btb_prediction_Freg_Tcu), .Z(n5)
         );
  Datapath_NBIT_DATA32_NBIT_IRAM_ADDR5 DP ( .DP_enable(DLX_enable), .DP_clk(
        DLX_clk), .DP_reset(DLX_reset), .DP_btb_target_prediction(
        s_target_prediction_Fbtb_Tdp), .DP_btb_prediction(
        s_btb_prediction_Fbtb_Treg), .DP_IR(DLX_IR), .DP_Rd1(
        s_DE_cw_Fcu_Tdp[1]), .DP_Rd2(s_DE_cw_Fcu_Tdp[2]), .DP_Wr(
        s_DE_cw_Fcu_Tdp[3]), .DP_JMP_branch(s_DE_cw_Fcu_Tdp[4:5]), 
        .DP_sign_extender(s_DE_cw_Fcu_Tdp[6:7]), .DP_save_PC(s_save_PC_Fcu_Tdp), .DP_Shift_Amount_sel({s_EX_cw_Fcu_Tdp[8], n7}), .DP_use_immediate(
        s_use_immediate_Fcu_Tdp), .DP_reverse_operands(n7), .DP_ALU_Opcode(
        s_EX_cw_Fcu_Tdp[10:15]), .DP_EX_enable(s_EX_cw_Fcu_Tdp[16]), 
        .DP_UUW_sel(s_MEM_cw_Fcu_Tdp), .DP_Store_reduce(s_MEM_cw_Fcu_Tdp_21), 
        .DP_Store_BYTE_half(s_MEM_cw_Fcu_Tdp_22), .DP_Load_data_from_DRAM(
        DLX_read_data), .DP_WB_sel(s_WB_cw_Fcu_Tdp[23]), .DP_Load_reduce(
        s_WB_cw_Fcu_Tdp[24]), .DP_Load_BYTE_half(s_WB_cw_Fcu_Tdp[25]), 
        .DP_Load_SGN_usg_reduce(s_WB_cw_Fcu_Tdp[26]), .DP_insert_bubble(
        s_insert_bubble_Fdp_Tcu), .DP_PC(DLX_PC), .DP_IF_ID_instr_is_branch(
        s_IFID_istr_is_brnch_Fdp_Tbmm), .DP_IR_opcode(s_IR_opcode_Fdp_Tcu), 
        .DP_IR_func(s_IR_func_Fdp_Tcu), .DP_restore_BTB(s_restore_Fdp_Tbmm), 
        .DP_branch_taken(s_branch_taken_Fdp_Tdp_cu), .DP_computed_new_PC(
        s_computed_NPC_Fdp_Tbmm), .DP_data_to_DRAM(DLX_written_data), 
        .DP_address_to_DRAM(DLX_address_written_data) );
  Reg1Bit_0 REG_BTB_PRED ( .clk(DLX_clk), .reset(n6), .data_in(
        s_btb_prediction_Fbtb_Treg), .enable(s_insert_bubble_Fdp_Tcu), .load(
        1'b1), .data_out(s_btb_prediction_Freg_Tcu) );
  ControlUnit CU ( .CU_instr_opcode(s_IR_opcode_Fdp_Tcu), .CU_instr_func(
        s_IR_func_Fdp_Tcu), .CU_enable(DLX_enable), .CU_reset(n6), .CU_clk(
        DLX_clk), .CU_flush(s_flush), .CU_bubble(s_insert_bubble_Fdp_Tcu), 
        .CU_CW_DE(s_DE_cw_Fcu_Tdp), .CU_CW_EX(s_EX_cw_Fcu_Tdp), .CU_CW_MEM({
        s_MEM_cw_Fcu_Tdp, DLX_RD_wr_DRAM, DLX_enable_DRAM, s_MEM_cw_Fcu_Tdp_21, 
        s_MEM_cw_Fcu_Tdp_22}), .CU_CW_WB(s_WB_cw_Fcu_Tdp), .CU_error(DLX_error) );
  NRegister_N32_0 PC_reg ( .clk(DLX_clk), .reset(n6), .data_in(DLX_PC), 
        .enable(s_insert_bubble_Fdp_Tcu), .load(1'b1), .data_out(
        s_NPC_Fdp_Tbmm) );
  BTB_misprediction_manager_NBIT_PC32 BMM ( .BMM_clk(DLX_clk), .BMM_reset(n6), 
        .BMM_enable(s_insert_bubble_Fdp_Tcu), .BMM_restore(s_restore_Fdp_Tbmm), 
        .BMM_PC(DLX_PC), .BMM_NPC(s_NPC_Fdp_Tbmm), .BMM_computed_PC(
        s_computed_NPC_Fdp_Tbmm), .BMM_is_branch(s_IFID_istr_is_brnch_Fdp_Tbmm), .BMM_branch_taken(s_branch_taken_Fdp_Tdp_cu), .BMM_PC_BTB(s_PC_Fbmm_Tbtb), 
        .BMM_NPC_BTB(s_NPC_Fbmm_Tbtb), .BMM_computed_PC_BTB(
        s_computed_NPC_Fbmm_Tbtb), .BMM_restore_BTB(s_restore_Fbmm_Tbtb), 
        .BMM_is_branch_BTB(s_IFID_istr_is_brnch_Fbmm_Tbtb), 
        .BMM_branch_taken_BTB(s_branch_taken_Fd_bmm_Tbtb) );
  BTB_N_ENTRY32_NBIT_ENTRY32_NBIT_TARGET32_NBIT_PREDICTION3 BTB_cache ( 
        .BTB_clk(DLX_clk), .BTB_rst(n6), .BTB_enable(s_insert_bubble_Fdp_Tcu), 
        .BTB_restore(s_restore_Fbmm_Tbtb), .BTB_PC_From_IF(s_PC_Fbmm_Tbtb), 
        .BTB_PC_From_DE(s_NPC_Fbmm_Tbtb), .BTB_target_From_DE(
        s_computed_NPC_Fbmm_Tbtb), .BTB_is_branch(
        s_IFID_istr_is_brnch_Fbmm_Tbtb), .BTB_branch_taken(
        s_branch_taken_Fd_bmm_Tbtb), .BTB_target_prediction(
        s_target_prediction_Fbtb_Tdp), .BTB_prediction(
        s_btb_prediction_Fbtb_Treg) );
  BUF_X2 U10 ( .A(s_EX_cw_Fcu_Tdp[9]), .Z(n7) );
  BUF_X1 U11 ( .A(DLX_reset), .Z(n6) );
  AND2_X1 U12 ( .A1(s_DE_cw_Fcu_Tdp[9]), .A2(s_DE_cw_Fcu_Tdp[8]), .ZN(
        s_save_PC_Fcu_Tdp) );
  INV_X1 U13 ( .A(s_DE_cw_Fcu_Tdp[2]), .ZN(s_use_immediate_Fcu_Tdp) );
endmodule

